module disp(
            input clk,
            input display_en,
			input neg_en,
            input [15:0] tmp,
            output reg[7:0] digit0,
            output reg[7:0] digit1,
			output reg[7:0] digit2,
			output reg[7:0] digit3
            );
//definition of 7-segment display with order: h(point),g,f,e,d,c,b,a
parameter EMPTY=8'b00000000;
parameter ZERO=8'b00111111;
parameter ONE=8'b00000110;
parameter TWO=8'b01011011;
parameter THREE=8'b01001111;
parameter FOUR=8'b01100110;
parameter FIVE=8'b01101101;
parameter SIX=8'b01111101;
parameter SEVEN=8'b00000111;
parameter EIGHT=8'b01111111;
parameter NINE=8'b01101111;
parameter MIN=8'b01000000;
parameter E=8'b01111001;
parameter R=8'b01110111;

always @(posedge clk)
begin
  if (display_en & ~neg_en)
    case (tmp)
      16'd10000:begin digit0<=R; digit1<=R; digit2<=E; digit3<=EMPTY; end
      16'd0: begin digit0<=ZERO; digit1<=EMPTY; digit2<=EMPTY; digit3<=EMPTY; end
      16'd1: begin digit0<=ONE; digit1<=EMPTY; digit2<=EMPTY; digit3<=EMPTY; end
      16'd2: begin digit0<=TWO; digit1<=EMPTY; digit2<=EMPTY; digit3<=EMPTY; end
      16'd3: begin digit0<=THREE; digit1<=EMPTY; digit2<=EMPTY; digit3<=EMPTY; end
      16'd4: begin digit0<=FOUR; digit1<=EMPTY; digit2<=EMPTY; digit3<=EMPTY; end
      16'd5: begin digit0<=FIVE; digit1<=EMPTY; digit2<=EMPTY; digit3<=EMPTY; end
      16'd6: begin digit0<=SIX; digit1<=EMPTY; digit2<=EMPTY; digit3<=EMPTY; end
      16'd7: begin digit0<=SEVEN; digit1<=EMPTY; digit2<=EMPTY; digit3<=EMPTY; end
      16'd8: begin digit0<=EIGHT; digit1<=EMPTY; digit2<=EMPTY; digit3<=EMPTY; end
      16'd9: begin digit0<=NINE; digit1<=EMPTY; digit2<=EMPTY; digit3<=EMPTY; end
      16'd10: begin digit0<=ZERO; digit1<=ONE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd11: begin digit0<=ONE; digit1<=ONE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd12: begin digit0<=TWO; digit1<=ONE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd13: begin digit0<=THREE; digit1<=ONE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd14: begin digit0<=FOUR; digit1<=ONE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd15: begin digit0<=FIVE; digit1<=ONE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd16: begin digit0<=SIX; digit1<=ONE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd17: begin digit0<=SEVEN; digit1<=ONE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd18: begin digit0<=EIGHT; digit1<=ONE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd19: begin digit0<=NINE; digit1<=ONE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd20: begin digit0<=ZERO; digit1<=TWO; digit2<=EMPTY; digit3<=EMPTY; end
      16'd21: begin digit0<=ONE; digit1<=TWO; digit2<=EMPTY; digit3<=EMPTY; end
      16'd22: begin digit0<=TWO; digit1<=TWO; digit2<=EMPTY; digit3<=EMPTY; end
      16'd23: begin digit0<=THREE; digit1<=TWO; digit2<=EMPTY; digit3<=EMPTY; end
      16'd24: begin digit0<=FOUR; digit1<=TWO; digit2<=EMPTY; digit3<=EMPTY; end
      16'd25: begin digit0<=FIVE; digit1<=TWO; digit2<=EMPTY; digit3<=EMPTY; end
      16'd26: begin digit0<=SIX; digit1<=TWO; digit2<=EMPTY; digit3<=EMPTY; end
      16'd27: begin digit0<=SEVEN; digit1<=TWO; digit2<=EMPTY; digit3<=EMPTY; end
      16'd28: begin digit0<=EIGHT; digit1<=TWO; digit2<=EMPTY; digit3<=EMPTY; end
      16'd29: begin digit0<=NINE; digit1<=TWO; digit2<=EMPTY; digit3<=EMPTY; end
      16'd30: begin digit0<=ZERO; digit1<=THREE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd31: begin digit0<=ONE; digit1<=THREE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd32: begin digit0<=TWO; digit1<=THREE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd33: begin digit0<=THREE; digit1<=THREE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd34: begin digit0<=FOUR; digit1<=THREE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd35: begin digit0<=FIVE; digit1<=THREE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd36: begin digit0<=SIX; digit1<=THREE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd37: begin digit0<=SEVEN; digit1<=THREE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd38: begin digit0<=EIGHT; digit1<=THREE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd39: begin digit0<=NINE; digit1<=THREE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd40: begin digit0<=ZERO; digit1<=FOUR; digit2<=EMPTY; digit3<=EMPTY; end
      16'd41: begin digit0<=ONE; digit1<=FOUR; digit2<=EMPTY; digit3<=EMPTY; end
      16'd42: begin digit0<=TWO; digit1<=FOUR; digit2<=EMPTY; digit3<=EMPTY; end
      16'd43: begin digit0<=THREE; digit1<=FOUR; digit2<=EMPTY; digit3<=EMPTY; end
      16'd44: begin digit0<=FOUR; digit1<=FOUR; digit2<=EMPTY; digit3<=EMPTY; end
      16'd45: begin digit0<=FIVE; digit1<=FOUR; digit2<=EMPTY; digit3<=EMPTY; end
      16'd46: begin digit0<=SIX; digit1<=FOUR; digit2<=EMPTY; digit3<=EMPTY; end
      16'd47: begin digit0<=SEVEN; digit1<=FOUR; digit2<=EMPTY; digit3<=EMPTY; end
      16'd48: begin digit0<=EIGHT; digit1<=FOUR; digit2<=EMPTY; digit3<=EMPTY; end
      16'd49: begin digit0<=NINE; digit1<=FOUR; digit2<=EMPTY; digit3<=EMPTY; end
      16'd50: begin digit0<=ZERO; digit1<=FIVE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd51: begin digit0<=ONE; digit1<=FIVE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd52: begin digit0<=TWO; digit1<=FIVE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd53: begin digit0<=THREE; digit1<=FIVE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd54: begin digit0<=FOUR; digit1<=FIVE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd55: begin digit0<=FIVE; digit1<=FIVE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd56: begin digit0<=SIX; digit1<=FIVE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd57: begin digit0<=SEVEN; digit1<=FIVE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd58: begin digit0<=EIGHT; digit1<=FIVE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd59: begin digit0<=NINE; digit1<=FIVE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd60: begin digit0<=ZERO; digit1<=SIX; digit2<=EMPTY; digit3<=EMPTY; end
      16'd61: begin digit0<=ONE; digit1<=SIX; digit2<=EMPTY; digit3<=EMPTY; end
      16'd62: begin digit0<=TWO; digit1<=SIX; digit2<=EMPTY; digit3<=EMPTY; end
      16'd63: begin digit0<=THREE; digit1<=SIX; digit2<=EMPTY; digit3<=EMPTY; end
      16'd64: begin digit0<=FOUR; digit1<=SIX; digit2<=EMPTY; digit3<=EMPTY; end
      16'd65: begin digit0<=FIVE; digit1<=SIX; digit2<=EMPTY; digit3<=EMPTY; end
      16'd66: begin digit0<=SIX; digit1<=SIX; digit2<=EMPTY; digit3<=EMPTY; end
      16'd67: begin digit0<=SEVEN; digit1<=SIX; digit2<=EMPTY; digit3<=EMPTY; end
      16'd68: begin digit0<=EIGHT; digit1<=SIX; digit2<=EMPTY; digit3<=EMPTY; end
      16'd69: begin digit0<=NINE; digit1<=SIX; digit2<=EMPTY; digit3<=EMPTY; end
      16'd70: begin digit0<=ZERO; digit1<=SEVEN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd71: begin digit0<=ONE; digit1<=SEVEN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd72: begin digit0<=TWO; digit1<=SEVEN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd73: begin digit0<=THREE; digit1<=SEVEN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd74: begin digit0<=FOUR; digit1<=SEVEN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd75: begin digit0<=FIVE; digit1<=SEVEN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd76: begin digit0<=SIX; digit1<=SEVEN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd77: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd78: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd79: begin digit0<=NINE; digit1<=SEVEN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd80: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EMPTY; digit3<=EMPTY; end
      16'd81: begin digit0<=ONE; digit1<=EIGHT; digit2<=EMPTY; digit3<=EMPTY; end
      16'd82: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EMPTY; digit3<=EMPTY; end
      16'd83: begin digit0<=THREE; digit1<=EIGHT; digit2<=EMPTY; digit3<=EMPTY; end
      16'd84: begin digit0<=FOUR; digit1<=EIGHT; digit2<=EMPTY; digit3<=EMPTY; end
      16'd85: begin digit0<=FIVE; digit1<=EIGHT; digit2<=EMPTY; digit3<=EMPTY; end
      16'd86: begin digit0<=SIX; digit1<=EIGHT; digit2<=EMPTY; digit3<=EMPTY; end
      16'd87: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=EMPTY; digit3<=EMPTY; end
      16'd88: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=EMPTY; digit3<=EMPTY; end
      16'd89: begin digit0<=NINE; digit1<=EIGHT; digit2<=EMPTY; digit3<=EMPTY; end
      16'd90: begin digit0<=ZERO; digit1<=NINE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd91: begin digit0<=ONE; digit1<=NINE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd92: begin digit0<=ZERO; digit1<=NINE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd93: begin digit0<=THREE; digit1<=NINE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd94: begin digit0<=FOUR; digit1<=NINE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd95: begin digit0<=FIVE; digit1<=NINE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd96: begin digit0<=SIX; digit1<=NINE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd97: begin digit0<=SEVEN; digit1<=NINE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd98: begin digit0<=EIGHT; digit1<=NINE; digit2<=EMPTY; digit3<=EMPTY; end
      16'd99: begin digit0<=NINE; digit1<=NINE; digit2<=EMPTY; digit3<=EMPTY; end
	  16'd100: begin digit0<=ZERO; digit1<=ZERO; digit2<=ONE; digit3<=EMPTY; end
      16'd101: begin digit0<=ONE; digit1<=ZERO; digit2<=ONE; digit3<=EMPTY; end
      16'd102: begin digit0<=TWO; digit1<=ZERO; digit2<=ONE; digit3<=EMPTY; end
      16'd103: begin digit0<=THREE; digit1<=ZERO; digit2<=ONE; digit3<=EMPTY; end
      16'd104: begin digit0<=FOUR; digit1<=ZERO; digit2<=ONE; digit3<=EMPTY; end
      16'd105: begin digit0<=FIVE; digit1<=ZERO; digit2<=ONE; digit3<=EMPTY; end
      16'd106: begin digit0<=SIX; digit1<=ZERO; digit2<=ONE; digit3<=EMPTY; end
      16'd107: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ONE; digit3<=EMPTY; end
      16'd108: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ONE; digit3<=EMPTY; end
      16'd109: begin digit0<=NINE; digit1<=ZERO; digit2<=ONE; digit3<=EMPTY; end
      16'd110: begin digit0<=ZERO; digit1<=ONE; digit2<=ONE; digit3<=EMPTY; end
      16'd111: begin digit0<=ONE; digit1<=ONE; digit2<=ONE; digit3<=EMPTY; end
      16'd112: begin digit0<=TWO; digit1<=ONE; digit2<=ONE; digit3<=EMPTY; end
      16'd113: begin digit0<=THREE; digit1<=ONE; digit2<=ONE; digit3<=EMPTY; end
      16'd114: begin digit0<=FOUR; digit1<=ONE; digit2<=ONE; digit3<=EMPTY; end
      16'd115: begin digit0<=FIVE; digit1<=ONE; digit2<=ONE; digit3<=EMPTY; end
      16'd116: begin digit0<=SIX; digit1<=ONE; digit2<=ONE; digit3<=EMPTY; end
      16'd117: begin digit0<=SEVEN; digit1<=ONE; digit2<=ONE; digit3<=EMPTY; end
      16'd118: begin digit0<=EIGHT; digit1<=ONE; digit2<=ONE; digit3<=EMPTY; end
      16'd119: begin digit0<=NINE; digit1<=ONE; digit2<=ONE; digit3<=EMPTY; end
      16'd120: begin digit0<=ZERO; digit1<=TWO; digit2<=ONE; digit3<=EMPTY; end
      16'd121: begin digit0<=ONE; digit1<=TWO; digit2<=ONE; digit3<=EMPTY; end
      16'd122: begin digit0<=TWO; digit1<=TWO; digit2<=ONE; digit3<=EMPTY; end
      16'd123: begin digit0<=THREE; digit1<=TWO; digit2<=ONE; digit3<=EMPTY; end
      16'd124: begin digit0<=FOUR; digit1<=TWO; digit2<=ONE; digit3<=EMPTY; end
      16'd125: begin digit0<=FIVE; digit1<=TWO; digit2<=ONE; digit3<=EMPTY; end
      16'd126: begin digit0<=SIX; digit1<=TWO; digit2<=ONE; digit3<=EMPTY; end
      16'd127: begin digit0<=SEVEN; digit1<=TWO; digit2<=ONE; digit3<=EMPTY; end
      16'd128: begin digit0<=EIGHT; digit1<=TWO; digit2<=ONE; digit3<=EMPTY; end
      16'd129: begin digit0<=NINE; digit1<=TWO; digit2<=ONE; digit3<=EMPTY; end
      16'd130: begin digit0<=ZERO; digit1<=THREE; digit2<=ONE; digit3<=EMPTY; end
      16'd131: begin digit0<=ONE; digit1<=THREE; digit2<=ONE; digit3<=EMPTY; end
      16'd132: begin digit0<=TWO; digit1<=THREE; digit2<=ONE; digit3<=EMPTY; end
      16'd133: begin digit0<=THREE; digit1<=THREE; digit2<=ONE; digit3<=EMPTY; end
      16'd134: begin digit0<=FOUR; digit1<=THREE; digit2<=ONE; digit3<=EMPTY; end
      16'd135: begin digit0<=FIVE; digit1<=THREE; digit2<=ONE; digit3<=EMPTY; end
      16'd136: begin digit0<=SIX; digit1<=THREE; digit2<=ONE; digit3<=EMPTY; end
      16'd137: begin digit0<=SEVEN; digit1<=THREE; digit2<=ONE; digit3<=EMPTY; end
      16'd138: begin digit0<=EIGHT; digit1<=THREE; digit2<=ONE; digit3<=EMPTY; end
      16'd139: begin digit0<=NINE; digit1<=THREE; digit2<=ONE; digit3<=EMPTY; end
      16'd140: begin digit0<=ZERO; digit1<=FOUR; digit2<=ONE; digit3<=EMPTY; end
      16'd141: begin digit0<=ONE; digit1<=FOUR; digit2<=ONE; digit3<=EMPTY; end
      16'd142: begin digit0<=TWO; digit1<=FOUR; digit2<=ONE; digit3<=EMPTY; end
      16'd143: begin digit0<=THREE; digit1<=FOUR; digit2<=ONE; digit3<=EMPTY; end
      16'd144: begin digit0<=FOUR; digit1<=FOUR; digit2<=ONE; digit3<=EMPTY; end
      16'd145: begin digit0<=FIVE; digit1<=FOUR; digit2<=ONE; digit3<=EMPTY; end
      16'd146: begin digit0<=SIX; digit1<=FOUR; digit2<=ONE; digit3<=EMPTY; end
      16'd147: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ONE; digit3<=EMPTY; end
      16'd148: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ONE; digit3<=EMPTY; end
      16'd149: begin digit0<=NINE; digit1<=FOUR; digit2<=ONE; digit3<=EMPTY; end
      16'd150: begin digit0<=ZERO; digit1<=FIVE; digit2<=ONE; digit3<=EMPTY; end
      16'd151: begin digit0<=ONE; digit1<=FIVE; digit2<=ONE; digit3<=EMPTY; end
      16'd152: begin digit0<=TWO; digit1<=FIVE; digit2<=ONE; digit3<=EMPTY; end
      16'd153: begin digit0<=THREE; digit1<=FIVE; digit2<=ONE; digit3<=EMPTY; end
      16'd154: begin digit0<=FOUR; digit1<=FIVE; digit2<=ONE; digit3<=EMPTY; end
      16'd155: begin digit0<=FIVE; digit1<=FIVE; digit2<=ONE; digit3<=EMPTY; end
      16'd156: begin digit0<=SIX; digit1<=FIVE; digit2<=ONE; digit3<=EMPTY; end
      16'd157: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ONE; digit3<=EMPTY; end
      16'd158: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ONE; digit3<=EMPTY; end
      16'd159: begin digit0<=NINE; digit1<=FIVE; digit2<=ONE; digit3<=EMPTY; end
      16'd160: begin digit0<=ZERO; digit1<=SIX; digit2<=ONE; digit3<=EMPTY; end
      16'd161: begin digit0<=ONE; digit1<=SIX; digit2<=ONE; digit3<=EMPTY; end
      16'd162: begin digit0<=TWO; digit1<=SIX; digit2<=ONE; digit3<=EMPTY; end
      16'd163: begin digit0<=THREE; digit1<=SIX; digit2<=ONE; digit3<=EMPTY; end
      16'd164: begin digit0<=FOUR; digit1<=SIX; digit2<=ONE; digit3<=EMPTY; end
      16'd165: begin digit0<=FIVE; digit1<=SIX; digit2<=ONE; digit3<=EMPTY; end
      16'd166: begin digit0<=SIX; digit1<=SIX; digit2<=ONE; digit3<=EMPTY; end
      16'd167: begin digit0<=SEVEN; digit1<=SIX; digit2<=ONE; digit3<=EMPTY; end
      16'd168: begin digit0<=EIGHT; digit1<=SIX; digit2<=ONE; digit3<=EMPTY; end
      16'd169: begin digit0<=NINE; digit1<=SIX; digit2<=ONE; digit3<=EMPTY; end
      16'd170: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ONE; digit3<=EMPTY; end
      16'd171: begin digit0<=ONE; digit1<=SEVEN; digit2<=ONE; digit3<=EMPTY; end
      16'd172: begin digit0<=TWO; digit1<=SEVEN; digit2<=ONE; digit3<=EMPTY; end
      16'd173: begin digit0<=THREE; digit1<=SEVEN; digit2<=ONE; digit3<=EMPTY; end
      16'd174: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ONE; digit3<=EMPTY; end
      16'd175: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ONE; digit3<=EMPTY; end
      16'd176: begin digit0<=SIX; digit1<=SEVEN; digit2<=ONE; digit3<=EMPTY; end
      16'd177: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ONE; digit3<=EMPTY; end
      16'd178: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ONE; digit3<=EMPTY; end
      16'd179: begin digit0<=NINE; digit1<=SEVEN; digit2<=ONE; digit3<=EMPTY; end
      16'd180: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=EMPTY; end
      16'd181: begin digit0<=ONE; digit1<=EIGHT; digit2<=ONE; digit3<=EMPTY; end
      16'd182: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=EMPTY; end
      16'd183: begin digit0<=THREE; digit1<=EIGHT; digit2<=ONE; digit3<=EMPTY; end
      16'd184: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ONE; digit3<=EMPTY; end
      16'd185: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ONE; digit3<=EMPTY; end
      16'd186: begin digit0<=SIX; digit1<=EIGHT; digit2<=ONE; digit3<=EMPTY; end
      16'd187: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ONE; digit3<=EMPTY; end
      16'd188: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ONE; digit3<=EMPTY; end
      16'd189: begin digit0<=NINE; digit1<=EIGHT; digit2<=ONE; digit3<=EMPTY; end
      16'd190: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=EMPTY; end
      16'd191: begin digit0<=ONE; digit1<=NINE; digit2<=ONE; digit3<=EMPTY; end
      16'd192: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=EMPTY; end
      16'd193: begin digit0<=THREE; digit1<=NINE; digit2<=ONE; digit3<=EMPTY; end
      16'd194: begin digit0<=FOUR; digit1<=NINE; digit2<=ONE; digit3<=EMPTY; end
      16'd195: begin digit0<=FIVE; digit1<=NINE; digit2<=ONE; digit3<=EMPTY; end
      16'd196: begin digit0<=SIX; digit1<=NINE; digit2<=ONE; digit3<=EMPTY; end
      16'd197: begin digit0<=SEVEN; digit1<=NINE; digit2<=ONE; digit3<=EMPTY; end
      16'd198: begin digit0<=EIGHT; digit1<=NINE; digit2<=ONE; digit3<=EMPTY; end
      16'd199: begin digit0<=NINE; digit1<=NINE; digit2<=ONE; digit3<=EMPTY; end
	  16'd200: begin digit0<=ZERO; digit1<=ZERO; digit2<=TWO; digit3<=EMPTY; end
      16'd201: begin digit0<=ONE; digit1<=ZERO; digit2<=TWO; digit3<=EMPTY; end
      16'd202: begin digit0<=TWO; digit1<=ZERO; digit2<=TWO; digit3<=EMPTY; end
      16'd203: begin digit0<=THREE; digit1<=ZERO; digit2<=TWO; digit3<=EMPTY; end
      16'd204: begin digit0<=FOUR; digit1<=ZERO; digit2<=TWO; digit3<=EMPTY; end
      16'd205: begin digit0<=FIVE; digit1<=ZERO; digit2<=TWO; digit3<=EMPTY; end
      16'd206: begin digit0<=SIX; digit1<=ZERO; digit2<=TWO; digit3<=EMPTY; end
      16'd207: begin digit0<=SEVEN; digit1<=ZERO; digit2<=TWO; digit3<=EMPTY; end
      16'd208: begin digit0<=EIGHT; digit1<=ZERO; digit2<=TWO; digit3<=EMPTY; end
      16'd209: begin digit0<=NINE; digit1<=ZERO; digit2<=TWO; digit3<=EMPTY; end
      16'd210: begin digit0<=ZERO; digit1<=ONE; digit2<=TWO; digit3<=EMPTY; end
      16'd211: begin digit0<=ONE; digit1<=ONE; digit2<=TWO; digit3<=EMPTY; end
      16'd212: begin digit0<=TWO; digit1<=ONE; digit2<=TWO; digit3<=EMPTY; end
      16'd213: begin digit0<=THREE; digit1<=ONE; digit2<=TWO; digit3<=EMPTY; end
      16'd214: begin digit0<=FOUR; digit1<=ONE; digit2<=TWO; digit3<=EMPTY; end
      16'd215: begin digit0<=FIVE; digit1<=ONE; digit2<=TWO; digit3<=EMPTY; end
      16'd216: begin digit0<=SIX; digit1<=ONE; digit2<=TWO; digit3<=EMPTY; end
      16'd217: begin digit0<=SEVEN; digit1<=ONE; digit2<=TWO; digit3<=EMPTY; end
      16'd218: begin digit0<=EIGHT; digit1<=ONE; digit2<=TWO; digit3<=EMPTY; end
      16'd219: begin digit0<=NINE; digit1<=ONE; digit2<=TWO; digit3<=EMPTY; end
      16'd220: begin digit0<=ZERO; digit1<=TWO; digit2<=TWO; digit3<=EMPTY; end
      16'd221: begin digit0<=ONE; digit1<=TWO; digit2<=TWO; digit3<=EMPTY; end
      16'd222: begin digit0<=TWO; digit1<=TWO; digit2<=TWO; digit3<=EMPTY; end
      16'd223: begin digit0<=THREE; digit1<=TWO; digit2<=TWO; digit3<=EMPTY; end
      16'd224: begin digit0<=FOUR; digit1<=TWO; digit2<=TWO; digit3<=EMPTY; end
      16'd225: begin digit0<=FIVE; digit1<=TWO; digit2<=TWO; digit3<=EMPTY; end
      16'd226: begin digit0<=SIX; digit1<=TWO; digit2<=TWO; digit3<=EMPTY; end
      16'd227: begin digit0<=SEVEN; digit1<=TWO; digit2<=TWO; digit3<=EMPTY; end
      16'd228: begin digit0<=EIGHT; digit1<=TWO; digit2<=TWO; digit3<=EMPTY; end
      16'd229: begin digit0<=NINE; digit1<=TWO; digit2<=TWO; digit3<=EMPTY; end
      16'd230: begin digit0<=ZERO; digit1<=THREE; digit2<=TWO; digit3<=EMPTY; end
      16'd231: begin digit0<=ONE; digit1<=THREE; digit2<=TWO; digit3<=EMPTY; end
      16'd232: begin digit0<=TWO; digit1<=THREE; digit2<=TWO; digit3<=EMPTY; end
      16'd233: begin digit0<=THREE; digit1<=THREE; digit2<=TWO; digit3<=EMPTY; end
      16'd234: begin digit0<=FOUR; digit1<=THREE; digit2<=TWO; digit3<=EMPTY; end
      16'd235: begin digit0<=FIVE; digit1<=THREE; digit2<=TWO; digit3<=EMPTY; end
      16'd236: begin digit0<=SIX; digit1<=THREE; digit2<=TWO; digit3<=EMPTY; end
      16'd237: begin digit0<=SEVEN; digit1<=THREE; digit2<=TWO; digit3<=EMPTY; end
      16'd238: begin digit0<=EIGHT; digit1<=THREE; digit2<=TWO; digit3<=EMPTY; end
      16'd239: begin digit0<=NINE; digit1<=THREE; digit2<=TWO; digit3<=EMPTY; end
      16'd240: begin digit0<=ZERO; digit1<=FOUR; digit2<=TWO; digit3<=EMPTY; end
      16'd241: begin digit0<=ONE; digit1<=FOUR; digit2<=TWO; digit3<=EMPTY; end
      16'd242: begin digit0<=TWO; digit1<=FOUR; digit2<=TWO; digit3<=EMPTY; end
      16'd243: begin digit0<=THREE; digit1<=FOUR; digit2<=TWO; digit3<=EMPTY; end
      16'd244: begin digit0<=FOUR; digit1<=FOUR; digit2<=TWO; digit3<=EMPTY; end
      16'd245: begin digit0<=FIVE; digit1<=FOUR; digit2<=TWO; digit3<=EMPTY; end
      16'd246: begin digit0<=SIX; digit1<=FOUR; digit2<=TWO; digit3<=EMPTY; end
      16'd247: begin digit0<=SEVEN; digit1<=FOUR; digit2<=TWO; digit3<=EMPTY; end
      16'd248: begin digit0<=EIGHT; digit1<=FOUR; digit2<=TWO; digit3<=EMPTY; end
      16'd249: begin digit0<=NINE; digit1<=FOUR; digit2<=TWO; digit3<=EMPTY; end
      16'd250: begin digit0<=ZERO; digit1<=FIVE; digit2<=TWO; digit3<=EMPTY; end
      16'd251: begin digit0<=ONE; digit1<=FIVE; digit2<=TWO; digit3<=EMPTY; end
      16'd252: begin digit0<=TWO; digit1<=FIVE; digit2<=TWO; digit3<=EMPTY; end
      16'd253: begin digit0<=THREE; digit1<=FIVE; digit2<=TWO; digit3<=EMPTY; end
      16'd254: begin digit0<=FOUR; digit1<=FIVE; digit2<=TWO; digit3<=EMPTY; end
      16'd255: begin digit0<=FIVE; digit1<=FIVE; digit2<=TWO; digit3<=EMPTY; end
      16'd256: begin digit0<=SIX; digit1<=FIVE; digit2<=TWO; digit3<=EMPTY; end
      16'd257: begin digit0<=SEVEN; digit1<=FIVE; digit2<=TWO; digit3<=EMPTY; end
      16'd258: begin digit0<=EIGHT; digit1<=FIVE; digit2<=TWO; digit3<=EMPTY; end
      16'd259: begin digit0<=NINE; digit1<=FIVE; digit2<=TWO; digit3<=EMPTY; end
      16'd260: begin digit0<=ZERO; digit1<=SIX; digit2<=TWO; digit3<=EMPTY; end
      16'd261: begin digit0<=ONE; digit1<=SIX; digit2<=TWO; digit3<=EMPTY; end
      16'd262: begin digit0<=TWO; digit1<=SIX; digit2<=TWO; digit3<=EMPTY; end
      16'd263: begin digit0<=THREE; digit1<=SIX; digit2<=TWO; digit3<=EMPTY; end
      16'd264: begin digit0<=FOUR; digit1<=SIX; digit2<=TWO; digit3<=EMPTY; end
      16'd265: begin digit0<=FIVE; digit1<=SIX; digit2<=TWO; digit3<=EMPTY; end
      16'd266: begin digit0<=SIX; digit1<=SIX; digit2<=TWO; digit3<=EMPTY; end
      16'd267: begin digit0<=SEVEN; digit1<=SIX; digit2<=TWO; digit3<=EMPTY; end
      16'd268: begin digit0<=EIGHT; digit1<=SIX; digit2<=TWO; digit3<=EMPTY; end
      16'd269: begin digit0<=NINE; digit1<=SIX; digit2<=TWO; digit3<=EMPTY; end
      16'd270: begin digit0<=ZERO; digit1<=SEVEN; digit2<=TWO; digit3<=EMPTY; end
      16'd271: begin digit0<=ONE; digit1<=SEVEN; digit2<=TWO; digit3<=EMPTY; end
      16'd272: begin digit0<=TWO; digit1<=SEVEN; digit2<=TWO; digit3<=EMPTY; end
      16'd273: begin digit0<=THREE; digit1<=SEVEN; digit2<=TWO; digit3<=EMPTY; end
      16'd274: begin digit0<=FOUR; digit1<=SEVEN; digit2<=TWO; digit3<=EMPTY; end
      16'd275: begin digit0<=FIVE; digit1<=SEVEN; digit2<=TWO; digit3<=EMPTY; end
      16'd276: begin digit0<=SIX; digit1<=SEVEN; digit2<=TWO; digit3<=EMPTY; end
      16'd277: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=TWO; digit3<=EMPTY; end
      16'd278: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=TWO; digit3<=EMPTY; end
      16'd279: begin digit0<=NINE; digit1<=SEVEN; digit2<=TWO; digit3<=EMPTY; end
      16'd280: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=EMPTY; end
      16'd281: begin digit0<=ONE; digit1<=EIGHT; digit2<=TWO; digit3<=EMPTY; end
      16'd282: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=EMPTY; end
      16'd283: begin digit0<=THREE; digit1<=EIGHT; digit2<=TWO; digit3<=EMPTY; end
      16'd284: begin digit0<=FOUR; digit1<=EIGHT; digit2<=TWO; digit3<=EMPTY; end
      16'd285: begin digit0<=FIVE; digit1<=EIGHT; digit2<=TWO; digit3<=EMPTY; end
      16'd286: begin digit0<=SIX; digit1<=EIGHT; digit2<=TWO; digit3<=EMPTY; end
      16'd287: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=TWO; digit3<=EMPTY; end
      16'd288: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=TWO; digit3<=EMPTY; end
      16'd289: begin digit0<=NINE; digit1<=EIGHT; digit2<=TWO; digit3<=EMPTY; end
      16'd290: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=EMPTY; end
      16'd291: begin digit0<=ONE; digit1<=NINE; digit2<=TWO; digit3<=EMPTY; end
      16'd292: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=EMPTY; end
      16'd293: begin digit0<=THREE; digit1<=NINE; digit2<=TWO; digit3<=EMPTY; end
      16'd294: begin digit0<=FOUR; digit1<=NINE; digit2<=TWO; digit3<=EMPTY; end
      16'd295: begin digit0<=FIVE; digit1<=NINE; digit2<=TWO; digit3<=EMPTY; end
      16'd296: begin digit0<=SIX; digit1<=NINE; digit2<=TWO; digit3<=EMPTY; end
      16'd297: begin digit0<=SEVEN; digit1<=NINE; digit2<=TWO; digit3<=EMPTY; end
      16'd298: begin digit0<=EIGHT; digit1<=NINE; digit2<=TWO; digit3<=EMPTY; end
      16'd299: begin digit0<=NINE; digit1<=NINE; digit2<=TWO; digit3<=EMPTY; end
	  16'd300: begin digit0<=ZERO; digit1<=ZERO; digit2<=THREE; digit3<=EMPTY; end
      16'd301: begin digit0<=ONE; digit1<=ZERO; digit2<=THREE; digit3<=EMPTY; end
      16'd302: begin digit0<=TWO; digit1<=ZERO; digit2<=THREE; digit3<=EMPTY; end
      16'd303: begin digit0<=THREE; digit1<=ZERO; digit2<=THREE; digit3<=EMPTY; end
      16'd304: begin digit0<=FOUR; digit1<=ZERO; digit2<=THREE; digit3<=EMPTY; end
      16'd305: begin digit0<=FIVE; digit1<=ZERO; digit2<=THREE; digit3<=EMPTY; end
      16'd306: begin digit0<=SIX; digit1<=ZERO; digit2<=THREE; digit3<=EMPTY; end
      16'd307: begin digit0<=SEVEN; digit1<=ZERO; digit2<=THREE; digit3<=EMPTY; end
      16'd308: begin digit0<=EIGHT; digit1<=ZERO; digit2<=THREE; digit3<=EMPTY; end
      16'd309: begin digit0<=NINE; digit1<=ZERO; digit2<=THREE; digit3<=EMPTY; end
      16'd310: begin digit0<=ZERO; digit1<=ONE; digit2<=THREE; digit3<=EMPTY; end
      16'd311: begin digit0<=ONE; digit1<=ONE; digit2<=THREE; digit3<=EMPTY; end
      16'd312: begin digit0<=TWO; digit1<=ONE; digit2<=THREE; digit3<=EMPTY; end
      16'd313: begin digit0<=THREE; digit1<=ONE; digit2<=THREE; digit3<=EMPTY; end
      16'd314: begin digit0<=FOUR; digit1<=ONE; digit2<=THREE; digit3<=EMPTY; end
      16'd315: begin digit0<=FIVE; digit1<=ONE; digit2<=THREE; digit3<=EMPTY; end
      16'd316: begin digit0<=SIX; digit1<=ONE; digit2<=THREE; digit3<=EMPTY; end
      16'd317: begin digit0<=SEVEN; digit1<=ONE; digit2<=THREE; digit3<=EMPTY; end
      16'd318: begin digit0<=EIGHT; digit1<=ONE; digit2<=THREE; digit3<=EMPTY; end
      16'd319: begin digit0<=NINE; digit1<=ONE; digit2<=THREE; digit3<=EMPTY; end
      16'd320: begin digit0<=ZERO; digit1<=TWO; digit2<=THREE; digit3<=EMPTY; end
      16'd321: begin digit0<=ONE; digit1<=TWO; digit2<=THREE; digit3<=EMPTY; end
      16'd322: begin digit0<=TWO; digit1<=TWO; digit2<=THREE; digit3<=EMPTY; end
      16'd323: begin digit0<=THREE; digit1<=TWO; digit2<=THREE; digit3<=EMPTY; end
      16'd324: begin digit0<=FOUR; digit1<=TWO; digit2<=THREE; digit3<=EMPTY; end
      16'd325: begin digit0<=FIVE; digit1<=TWO; digit2<=THREE; digit3<=EMPTY; end
      16'd326: begin digit0<=SIX; digit1<=TWO; digit2<=THREE; digit3<=EMPTY; end
      16'd327: begin digit0<=SEVEN; digit1<=TWO; digit2<=THREE; digit3<=EMPTY; end
      16'd328: begin digit0<=EIGHT; digit1<=TWO; digit2<=THREE; digit3<=EMPTY; end
      16'd329: begin digit0<=NINE; digit1<=TWO; digit2<=THREE; digit3<=EMPTY; end
      16'd330: begin digit0<=ZERO; digit1<=THREE; digit2<=THREE; digit3<=EMPTY; end
      16'd331: begin digit0<=ONE; digit1<=THREE; digit2<=THREE; digit3<=EMPTY; end
      16'd332: begin digit0<=TWO; digit1<=THREE; digit2<=THREE; digit3<=EMPTY; end
      16'd333: begin digit0<=THREE; digit1<=THREE; digit2<=THREE; digit3<=EMPTY; end
      16'd334: begin digit0<=FOUR; digit1<=THREE; digit2<=THREE; digit3<=EMPTY; end
      16'd335: begin digit0<=FIVE; digit1<=THREE; digit2<=THREE; digit3<=EMPTY; end
      16'd336: begin digit0<=SIX; digit1<=THREE; digit2<=THREE; digit3<=EMPTY; end
      16'd337: begin digit0<=SEVEN; digit1<=THREE; digit2<=THREE; digit3<=EMPTY; end
      16'd338: begin digit0<=EIGHT; digit1<=THREE; digit2<=THREE; digit3<=EMPTY; end
      16'd339: begin digit0<=NINE; digit1<=THREE; digit2<=THREE; digit3<=EMPTY; end
      16'd340: begin digit0<=ZERO; digit1<=FOUR; digit2<=THREE; digit3<=EMPTY; end
      16'd341: begin digit0<=ONE; digit1<=FOUR; digit2<=THREE; digit3<=EMPTY; end
      16'd342: begin digit0<=TWO; digit1<=FOUR; digit2<=THREE; digit3<=EMPTY; end
      16'd343: begin digit0<=THREE; digit1<=FOUR; digit2<=THREE; digit3<=EMPTY; end
      16'd344: begin digit0<=FOUR; digit1<=FOUR; digit2<=THREE; digit3<=EMPTY; end
      16'd345: begin digit0<=FIVE; digit1<=FOUR; digit2<=THREE; digit3<=EMPTY; end
      16'd346: begin digit0<=SIX; digit1<=FOUR; digit2<=THREE; digit3<=EMPTY; end
      16'd347: begin digit0<=SEVEN; digit1<=FOUR; digit2<=THREE; digit3<=EMPTY; end
      16'd348: begin digit0<=EIGHT; digit1<=FOUR; digit2<=THREE; digit3<=EMPTY; end
      16'd349: begin digit0<=NINE; digit1<=FOUR; digit2<=THREE; digit3<=EMPTY; end
      16'd350: begin digit0<=ZERO; digit1<=FIVE; digit2<=THREE; digit3<=EMPTY; end
      16'd351: begin digit0<=ONE; digit1<=FIVE; digit2<=THREE; digit3<=EMPTY; end
      16'd352: begin digit0<=TWO; digit1<=FIVE; digit2<=THREE; digit3<=EMPTY; end
      16'd353: begin digit0<=THREE; digit1<=FIVE; digit2<=THREE; digit3<=EMPTY; end
      16'd354: begin digit0<=FOUR; digit1<=FIVE; digit2<=THREE; digit3<=EMPTY; end
      16'd355: begin digit0<=FIVE; digit1<=FIVE; digit2<=THREE; digit3<=EMPTY; end
      16'd356: begin digit0<=SIX; digit1<=FIVE; digit2<=THREE; digit3<=EMPTY; end
      16'd357: begin digit0<=SEVEN; digit1<=FIVE; digit2<=THREE; digit3<=EMPTY; end
      16'd358: begin digit0<=EIGHT; digit1<=FIVE; digit2<=THREE; digit3<=EMPTY; end
      16'd359: begin digit0<=NINE; digit1<=FIVE; digit2<=THREE; digit3<=EMPTY; end
      16'd360: begin digit0<=ZERO; digit1<=SIX; digit2<=THREE; digit3<=EMPTY; end
      16'd361: begin digit0<=ONE; digit1<=SIX; digit2<=THREE; digit3<=EMPTY; end
      16'd362: begin digit0<=TWO; digit1<=SIX; digit2<=THREE; digit3<=EMPTY; end
      16'd363: begin digit0<=THREE; digit1<=SIX; digit2<=THREE; digit3<=EMPTY; end
      16'd364: begin digit0<=FOUR; digit1<=SIX; digit2<=THREE; digit3<=EMPTY; end
      16'd365: begin digit0<=FIVE; digit1<=SIX; digit2<=THREE; digit3<=EMPTY; end
      16'd366: begin digit0<=SIX; digit1<=SIX; digit2<=THREE; digit3<=EMPTY; end
      16'd367: begin digit0<=SEVEN; digit1<=SIX; digit2<=THREE; digit3<=EMPTY; end
      16'd368: begin digit0<=EIGHT; digit1<=SIX; digit2<=THREE; digit3<=EMPTY; end
      16'd369: begin digit0<=NINE; digit1<=SIX; digit2<=THREE; digit3<=EMPTY; end
      16'd370: begin digit0<=ZERO; digit1<=SEVEN; digit2<=THREE; digit3<=EMPTY; end
      16'd371: begin digit0<=ONE; digit1<=SEVEN; digit2<=THREE; digit3<=EMPTY; end
      16'd372: begin digit0<=TWO; digit1<=SEVEN; digit2<=THREE; digit3<=EMPTY; end
      16'd373: begin digit0<=THREE; digit1<=SEVEN; digit2<=THREE; digit3<=EMPTY; end
      16'd374: begin digit0<=FOUR; digit1<=SEVEN; digit2<=THREE; digit3<=EMPTY; end
      16'd375: begin digit0<=FIVE; digit1<=SEVEN; digit2<=THREE; digit3<=EMPTY; end
      16'd376: begin digit0<=SIX; digit1<=SEVEN; digit2<=THREE; digit3<=EMPTY; end
      16'd377: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=THREE; digit3<=EMPTY; end
      16'd378: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=THREE; digit3<=EMPTY; end
      16'd379: begin digit0<=NINE; digit1<=SEVEN; digit2<=THREE; digit3<=EMPTY; end
      16'd380: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=EMPTY; end
      16'd381: begin digit0<=ONE; digit1<=EIGHT; digit2<=THREE; digit3<=EMPTY; end
      16'd382: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=EMPTY; end
      16'd383: begin digit0<=THREE; digit1<=EIGHT; digit2<=THREE; digit3<=EMPTY; end
      16'd384: begin digit0<=FOUR; digit1<=EIGHT; digit2<=THREE; digit3<=EMPTY; end
      16'd385: begin digit0<=FIVE; digit1<=EIGHT; digit2<=THREE; digit3<=EMPTY; end
      16'd386: begin digit0<=SIX; digit1<=EIGHT; digit2<=THREE; digit3<=EMPTY; end
      16'd387: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=THREE; digit3<=EMPTY; end
      16'd388: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=THREE; digit3<=EMPTY; end
      16'd389: begin digit0<=NINE; digit1<=EIGHT; digit2<=THREE; digit3<=EMPTY; end
      16'd390: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=EMPTY; end
      16'd391: begin digit0<=ONE; digit1<=NINE; digit2<=THREE; digit3<=EMPTY; end
      16'd392: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=EMPTY; end
      16'd393: begin digit0<=THREE; digit1<=NINE; digit2<=THREE; digit3<=EMPTY; end
      16'd394: begin digit0<=FOUR; digit1<=NINE; digit2<=THREE; digit3<=EMPTY; end
      16'd395: begin digit0<=FIVE; digit1<=NINE; digit2<=THREE; digit3<=EMPTY; end
      16'd396: begin digit0<=SIX; digit1<=NINE; digit2<=THREE; digit3<=EMPTY; end
      16'd397: begin digit0<=SEVEN; digit1<=NINE; digit2<=THREE; digit3<=EMPTY; end
      16'd398: begin digit0<=EIGHT; digit1<=NINE; digit2<=THREE; digit3<=EMPTY; end
      16'd399: begin digit0<=NINE; digit1<=NINE; digit2<=THREE; digit3<=EMPTY; end
	  16'd400: begin digit0<=ZERO; digit1<=ZERO; digit2<=FOUR; digit3<=EMPTY; end
      16'd401: begin digit0<=ONE; digit1<=ZERO; digit2<=FOUR; digit3<=EMPTY; end
      16'd402: begin digit0<=TWO; digit1<=ZERO; digit2<=FOUR; digit3<=EMPTY; end
      16'd403: begin digit0<=THREE; digit1<=ZERO; digit2<=FOUR; digit3<=EMPTY; end
      16'd404: begin digit0<=FOUR; digit1<=ZERO; digit2<=FOUR; digit3<=EMPTY; end
      16'd405: begin digit0<=FIVE; digit1<=ZERO; digit2<=FOUR; digit3<=EMPTY; end
      16'd406: begin digit0<=SIX; digit1<=ZERO; digit2<=FOUR; digit3<=EMPTY; end
      16'd407: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FOUR; digit3<=EMPTY; end
      16'd408: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FOUR; digit3<=EMPTY; end
      16'd409: begin digit0<=NINE; digit1<=ZERO; digit2<=FOUR; digit3<=EMPTY; end
      16'd410: begin digit0<=ZERO; digit1<=ONE; digit2<=FOUR; digit3<=EMPTY; end
      16'd411: begin digit0<=ONE; digit1<=ONE; digit2<=FOUR; digit3<=EMPTY; end
      16'd412: begin digit0<=TWO; digit1<=ONE; digit2<=FOUR; digit3<=EMPTY; end
      16'd413: begin digit0<=THREE; digit1<=ONE; digit2<=FOUR; digit3<=EMPTY; end
      16'd414: begin digit0<=FOUR; digit1<=ONE; digit2<=FOUR; digit3<=EMPTY; end
      16'd415: begin digit0<=FIVE; digit1<=ONE; digit2<=FOUR; digit3<=EMPTY; end
      16'd416: begin digit0<=SIX; digit1<=ONE; digit2<=FOUR; digit3<=EMPTY; end
      16'd417: begin digit0<=SEVEN; digit1<=ONE; digit2<=FOUR; digit3<=EMPTY; end
      16'd418: begin digit0<=EIGHT; digit1<=ONE; digit2<=FOUR; digit3<=EMPTY; end
      16'd419: begin digit0<=NINE; digit1<=ONE; digit2<=FOUR; digit3<=EMPTY; end
      16'd420: begin digit0<=ZERO; digit1<=TWO; digit2<=FOUR; digit3<=EMPTY; end
      16'd421: begin digit0<=ONE; digit1<=TWO; digit2<=FOUR; digit3<=EMPTY; end
      16'd422: begin digit0<=TWO; digit1<=TWO; digit2<=FOUR; digit3<=EMPTY; end
      16'd423: begin digit0<=THREE; digit1<=TWO; digit2<=FOUR; digit3<=EMPTY; end
      16'd424: begin digit0<=FOUR; digit1<=TWO; digit2<=FOUR; digit3<=EMPTY; end
      16'd425: begin digit0<=FIVE; digit1<=TWO; digit2<=FOUR; digit3<=EMPTY; end
      16'd426: begin digit0<=SIX; digit1<=TWO; digit2<=FOUR; digit3<=EMPTY; end
      16'd427: begin digit0<=SEVEN; digit1<=TWO; digit2<=FOUR; digit3<=EMPTY; end
      16'd428: begin digit0<=EIGHT; digit1<=TWO; digit2<=FOUR; digit3<=EMPTY; end
      16'd429: begin digit0<=NINE; digit1<=TWO; digit2<=FOUR; digit3<=EMPTY; end
      16'd430: begin digit0<=ZERO; digit1<=THREE; digit2<=FOUR; digit3<=EMPTY; end
      16'd431: begin digit0<=ONE; digit1<=THREE; digit2<=FOUR; digit3<=EMPTY; end
      16'd432: begin digit0<=TWO; digit1<=THREE; digit2<=FOUR; digit3<=EMPTY; end
      16'd433: begin digit0<=THREE; digit1<=THREE; digit2<=FOUR; digit3<=EMPTY; end
      16'd434: begin digit0<=FOUR; digit1<=THREE; digit2<=FOUR; digit3<=EMPTY; end
      16'd435: begin digit0<=FIVE; digit1<=THREE; digit2<=FOUR; digit3<=EMPTY; end
      16'd436: begin digit0<=SIX; digit1<=THREE; digit2<=FOUR; digit3<=EMPTY; end
      16'd437: begin digit0<=SEVEN; digit1<=THREE; digit2<=FOUR; digit3<=EMPTY; end
      16'd438: begin digit0<=EIGHT; digit1<=THREE; digit2<=FOUR; digit3<=EMPTY; end
      16'd439: begin digit0<=NINE; digit1<=THREE; digit2<=FOUR; digit3<=EMPTY; end
      16'd440: begin digit0<=ZERO; digit1<=FOUR; digit2<=FOUR; digit3<=EMPTY; end
      16'd441: begin digit0<=ONE; digit1<=FOUR; digit2<=FOUR; digit3<=EMPTY; end
      16'd442: begin digit0<=TWO; digit1<=FOUR; digit2<=FOUR; digit3<=EMPTY; end
      16'd443: begin digit0<=THREE; digit1<=FOUR; digit2<=FOUR; digit3<=EMPTY; end
      16'd444: begin digit0<=FOUR; digit1<=FOUR; digit2<=FOUR; digit3<=EMPTY; end
      16'd445: begin digit0<=FIVE; digit1<=FOUR; digit2<=FOUR; digit3<=EMPTY; end
      16'd446: begin digit0<=SIX; digit1<=FOUR; digit2<=FOUR; digit3<=EMPTY; end
      16'd447: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FOUR; digit3<=EMPTY; end
      16'd448: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FOUR; digit3<=EMPTY; end
      16'd449: begin digit0<=NINE; digit1<=FOUR; digit2<=FOUR; digit3<=EMPTY; end
      16'd450: begin digit0<=ZERO; digit1<=FIVE; digit2<=FOUR; digit3<=EMPTY; end
      16'd451: begin digit0<=ONE; digit1<=FIVE; digit2<=FOUR; digit3<=EMPTY; end
      16'd452: begin digit0<=TWO; digit1<=FIVE; digit2<=FOUR; digit3<=EMPTY; end
      16'd453: begin digit0<=THREE; digit1<=FIVE; digit2<=FOUR; digit3<=EMPTY; end
      16'd454: begin digit0<=FOUR; digit1<=FIVE; digit2<=FOUR; digit3<=EMPTY; end
      16'd455: begin digit0<=FIVE; digit1<=FIVE; digit2<=FOUR; digit3<=EMPTY; end
      16'd456: begin digit0<=SIX; digit1<=FIVE; digit2<=FOUR; digit3<=EMPTY; end
      16'd457: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FOUR; digit3<=EMPTY; end
      16'd458: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FOUR; digit3<=EMPTY; end
      16'd459: begin digit0<=NINE; digit1<=FIVE; digit2<=FOUR; digit3<=EMPTY; end
      16'd460: begin digit0<=ZERO; digit1<=SIX; digit2<=FOUR; digit3<=EMPTY; end
      16'd461: begin digit0<=ONE; digit1<=SIX; digit2<=FOUR; digit3<=EMPTY; end
      16'd462: begin digit0<=TWO; digit1<=SIX; digit2<=FOUR; digit3<=EMPTY; end
      16'd463: begin digit0<=THREE; digit1<=SIX; digit2<=FOUR; digit3<=EMPTY; end
      16'd464: begin digit0<=FOUR; digit1<=SIX; digit2<=FOUR; digit3<=EMPTY; end
      16'd465: begin digit0<=FIVE; digit1<=SIX; digit2<=FOUR; digit3<=EMPTY; end
      16'd466: begin digit0<=SIX; digit1<=SIX; digit2<=FOUR; digit3<=EMPTY; end
      16'd467: begin digit0<=SEVEN; digit1<=SIX; digit2<=FOUR; digit3<=EMPTY; end
      16'd468: begin digit0<=EIGHT; digit1<=SIX; digit2<=FOUR; digit3<=EMPTY; end
      16'd469: begin digit0<=NINE; digit1<=SIX; digit2<=FOUR; digit3<=EMPTY; end
      16'd470: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FOUR; digit3<=EMPTY; end
      16'd471: begin digit0<=ONE; digit1<=SEVEN; digit2<=FOUR; digit3<=EMPTY; end
      16'd472: begin digit0<=TWO; digit1<=SEVEN; digit2<=FOUR; digit3<=EMPTY; end
      16'd473: begin digit0<=THREE; digit1<=SEVEN; digit2<=FOUR; digit3<=EMPTY; end
      16'd474: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FOUR; digit3<=EMPTY; end
      16'd475: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FOUR; digit3<=EMPTY; end
      16'd476: begin digit0<=SIX; digit1<=SEVEN; digit2<=FOUR; digit3<=EMPTY; end
      16'd477: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FOUR; digit3<=EMPTY; end
      16'd478: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FOUR; digit3<=EMPTY; end
      16'd479: begin digit0<=NINE; digit1<=SEVEN; digit2<=FOUR; digit3<=EMPTY; end
      16'd480: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=EMPTY; end
      16'd481: begin digit0<=ONE; digit1<=EIGHT; digit2<=FOUR; digit3<=EMPTY; end
      16'd482: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=EMPTY; end
      16'd483: begin digit0<=THREE; digit1<=EIGHT; digit2<=FOUR; digit3<=EMPTY; end
      16'd484: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FOUR; digit3<=EMPTY; end
      16'd485: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FOUR; digit3<=EMPTY; end
      16'd486: begin digit0<=SIX; digit1<=EIGHT; digit2<=FOUR; digit3<=EMPTY; end
      16'd487: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FOUR; digit3<=EMPTY; end
      16'd488: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FOUR; digit3<=EMPTY; end
      16'd489: begin digit0<=NINE; digit1<=EIGHT; digit2<=FOUR; digit3<=EMPTY; end
      16'd490: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=EMPTY; end
      16'd491: begin digit0<=ONE; digit1<=NINE; digit2<=FOUR; digit3<=EMPTY; end
      16'd492: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=EMPTY; end
      16'd493: begin digit0<=THREE; digit1<=NINE; digit2<=FOUR; digit3<=EMPTY; end
      16'd494: begin digit0<=FOUR; digit1<=NINE; digit2<=FOUR; digit3<=EMPTY; end
      16'd495: begin digit0<=FIVE; digit1<=NINE; digit2<=FOUR; digit3<=EMPTY; end
      16'd496: begin digit0<=SIX; digit1<=NINE; digit2<=FOUR; digit3<=EMPTY; end
      16'd497: begin digit0<=SEVEN; digit1<=NINE; digit2<=FOUR; digit3<=EMPTY; end
      16'd498: begin digit0<=EIGHT; digit1<=NINE; digit2<=FOUR; digit3<=EMPTY; end
      16'd499: begin digit0<=NINE; digit1<=NINE; digit2<=FOUR; digit3<=EMPTY; end
	  16'd500: begin digit0<=ZERO; digit1<=ZERO; digit2<=FIVE; digit3<=EMPTY; end
      16'd501: begin digit0<=ONE; digit1<=ZERO; digit2<=FIVE; digit3<=EMPTY; end
      16'd502: begin digit0<=TWO; digit1<=ZERO; digit2<=FIVE; digit3<=EMPTY; end
      16'd503: begin digit0<=THREE; digit1<=ZERO; digit2<=FIVE; digit3<=EMPTY; end
      16'd504: begin digit0<=FOUR; digit1<=ZERO; digit2<=FIVE; digit3<=EMPTY; end
      16'd505: begin digit0<=FIVE; digit1<=ZERO; digit2<=FIVE; digit3<=EMPTY; end
      16'd506: begin digit0<=SIX; digit1<=ZERO; digit2<=FIVE; digit3<=EMPTY; end
      16'd507: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FIVE; digit3<=EMPTY; end
      16'd508: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FIVE; digit3<=EMPTY; end
      16'd509: begin digit0<=NINE; digit1<=ZERO; digit2<=FIVE; digit3<=EMPTY; end
      16'd510: begin digit0<=ZERO; digit1<=ONE; digit2<=FIVE; digit3<=EMPTY; end
      16'd511: begin digit0<=ONE; digit1<=ONE; digit2<=FIVE; digit3<=EMPTY; end
      16'd512: begin digit0<=TWO; digit1<=ONE; digit2<=FIVE; digit3<=EMPTY; end
      16'd513: begin digit0<=THREE; digit1<=ONE; digit2<=FIVE; digit3<=EMPTY; end
      16'd514: begin digit0<=FOUR; digit1<=ONE; digit2<=FIVE; digit3<=EMPTY; end
      16'd515: begin digit0<=FIVE; digit1<=ONE; digit2<=FIVE; digit3<=EMPTY; end
      16'd516: begin digit0<=SIX; digit1<=ONE; digit2<=FIVE; digit3<=EMPTY; end
      16'd517: begin digit0<=SEVEN; digit1<=ONE; digit2<=FIVE; digit3<=EMPTY; end
      16'd518: begin digit0<=EIGHT; digit1<=ONE; digit2<=FIVE; digit3<=EMPTY; end
      16'd519: begin digit0<=NINE; digit1<=ONE; digit2<=FIVE; digit3<=EMPTY; end
      16'd520: begin digit0<=ZERO; digit1<=TWO; digit2<=FIVE; digit3<=EMPTY; end
      16'd521: begin digit0<=ONE; digit1<=TWO; digit2<=FIVE; digit3<=EMPTY; end
      16'd522: begin digit0<=TWO; digit1<=TWO; digit2<=FIVE; digit3<=EMPTY; end
      16'd523: begin digit0<=THREE; digit1<=TWO; digit2<=FIVE; digit3<=EMPTY; end
      16'd524: begin digit0<=FOUR; digit1<=TWO; digit2<=FIVE; digit3<=EMPTY; end
      16'd525: begin digit0<=FIVE; digit1<=TWO; digit2<=FIVE; digit3<=EMPTY; end
      16'd526: begin digit0<=SIX; digit1<=TWO; digit2<=FIVE; digit3<=EMPTY; end
      16'd527: begin digit0<=SEVEN; digit1<=TWO; digit2<=FIVE; digit3<=EMPTY; end
      16'd528: begin digit0<=EIGHT; digit1<=TWO; digit2<=FIVE; digit3<=EMPTY; end
      16'd529: begin digit0<=NINE; digit1<=TWO; digit2<=FIVE; digit3<=EMPTY; end
      16'd530: begin digit0<=ZERO; digit1<=THREE; digit2<=FIVE; digit3<=EMPTY; end
      16'd531: begin digit0<=ONE; digit1<=THREE; digit2<=FIVE; digit3<=EMPTY; end
      16'd532: begin digit0<=TWO; digit1<=THREE; digit2<=FIVE; digit3<=EMPTY; end
      16'd533: begin digit0<=THREE; digit1<=THREE; digit2<=FIVE; digit3<=EMPTY; end
      16'd534: begin digit0<=FOUR; digit1<=THREE; digit2<=FIVE; digit3<=EMPTY; end
      16'd535: begin digit0<=FIVE; digit1<=THREE; digit2<=FIVE; digit3<=EMPTY; end
      16'd536: begin digit0<=SIX; digit1<=THREE; digit2<=FIVE; digit3<=EMPTY; end
      16'd537: begin digit0<=SEVEN; digit1<=THREE; digit2<=FIVE; digit3<=EMPTY; end
      16'd538: begin digit0<=EIGHT; digit1<=THREE; digit2<=FIVE; digit3<=EMPTY; end
      16'd539: begin digit0<=NINE; digit1<=THREE; digit2<=FIVE; digit3<=EMPTY; end
      16'd540: begin digit0<=ZERO; digit1<=FOUR; digit2<=FIVE; digit3<=EMPTY; end
      16'd541: begin digit0<=ONE; digit1<=FOUR; digit2<=FIVE; digit3<=EMPTY; end
      16'd542: begin digit0<=TWO; digit1<=FOUR; digit2<=FIVE; digit3<=EMPTY; end
      16'd543: begin digit0<=THREE; digit1<=FOUR; digit2<=FIVE; digit3<=EMPTY; end
      16'd544: begin digit0<=FOUR; digit1<=FOUR; digit2<=FIVE; digit3<=EMPTY; end
      16'd545: begin digit0<=FIVE; digit1<=FOUR; digit2<=FIVE; digit3<=EMPTY; end
      16'd546: begin digit0<=SIX; digit1<=FOUR; digit2<=FIVE; digit3<=EMPTY; end
      16'd547: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FIVE; digit3<=EMPTY; end
      16'd548: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FIVE; digit3<=EMPTY; end
      16'd549: begin digit0<=NINE; digit1<=FOUR; digit2<=FIVE; digit3<=EMPTY; end
      16'd550: begin digit0<=ZERO; digit1<=FIVE; digit2<=FIVE; digit3<=EMPTY; end
      16'd551: begin digit0<=ONE; digit1<=FIVE; digit2<=FIVE; digit3<=EMPTY; end
      16'd552: begin digit0<=TWO; digit1<=FIVE; digit2<=FIVE; digit3<=EMPTY; end
      16'd553: begin digit0<=THREE; digit1<=FIVE; digit2<=FIVE; digit3<=EMPTY; end
      16'd554: begin digit0<=FOUR; digit1<=FIVE; digit2<=FIVE; digit3<=EMPTY; end
      16'd555: begin digit0<=FIVE; digit1<=FIVE; digit2<=FIVE; digit3<=EMPTY; end
      16'd556: begin digit0<=SIX; digit1<=FIVE; digit2<=FIVE; digit3<=EMPTY; end
      16'd557: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FIVE; digit3<=EMPTY; end
      16'd558: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FIVE; digit3<=EMPTY; end
      16'd559: begin digit0<=NINE; digit1<=FIVE; digit2<=FIVE; digit3<=EMPTY; end
      16'd560: begin digit0<=ZERO; digit1<=SIX; digit2<=FIVE; digit3<=EMPTY; end
      16'd561: begin digit0<=ONE; digit1<=SIX; digit2<=FIVE; digit3<=EMPTY; end
      16'd562: begin digit0<=TWO; digit1<=SIX; digit2<=FIVE; digit3<=EMPTY; end
      16'd563: begin digit0<=THREE; digit1<=SIX; digit2<=FIVE; digit3<=EMPTY; end
      16'd564: begin digit0<=FOUR; digit1<=SIX; digit2<=FIVE; digit3<=EMPTY; end
      16'd565: begin digit0<=FIVE; digit1<=SIX; digit2<=FIVE; digit3<=EMPTY; end
      16'd566: begin digit0<=SIX; digit1<=SIX; digit2<=FIVE; digit3<=EMPTY; end
      16'd567: begin digit0<=SEVEN; digit1<=SIX; digit2<=FIVE; digit3<=EMPTY; end
      16'd568: begin digit0<=EIGHT; digit1<=SIX; digit2<=FIVE; digit3<=EMPTY; end
      16'd569: begin digit0<=NINE; digit1<=SIX; digit2<=FIVE; digit3<=EMPTY; end
      16'd570: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FIVE; digit3<=EMPTY; end
      16'd571: begin digit0<=ONE; digit1<=SEVEN; digit2<=FIVE; digit3<=EMPTY; end
      16'd572: begin digit0<=TWO; digit1<=SEVEN; digit2<=FIVE; digit3<=EMPTY; end
      16'd573: begin digit0<=THREE; digit1<=SEVEN; digit2<=FIVE; digit3<=EMPTY; end
      16'd574: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FIVE; digit3<=EMPTY; end
      16'd575: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FIVE; digit3<=EMPTY; end
      16'd576: begin digit0<=SIX; digit1<=SEVEN; digit2<=FIVE; digit3<=EMPTY; end
      16'd577: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FIVE; digit3<=EMPTY; end
      16'd578: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FIVE; digit3<=EMPTY; end
      16'd579: begin digit0<=NINE; digit1<=SEVEN; digit2<=FIVE; digit3<=EMPTY; end
      16'd580: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=EMPTY; end
      16'd581: begin digit0<=ONE; digit1<=EIGHT; digit2<=FIVE; digit3<=EMPTY; end
      16'd582: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=EMPTY; end
      16'd583: begin digit0<=THREE; digit1<=EIGHT; digit2<=FIVE; digit3<=EMPTY; end
      16'd584: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FIVE; digit3<=EMPTY; end
      16'd585: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FIVE; digit3<=EMPTY; end
      16'd586: begin digit0<=SIX; digit1<=EIGHT; digit2<=FIVE; digit3<=EMPTY; end
      16'd587: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FIVE; digit3<=EMPTY; end
      16'd588: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FIVE; digit3<=EMPTY; end
      16'd589: begin digit0<=NINE; digit1<=EIGHT; digit2<=FIVE; digit3<=EMPTY; end
      16'd590: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=EMPTY; end
      16'd591: begin digit0<=ONE; digit1<=NINE; digit2<=FIVE; digit3<=EMPTY; end
      16'd592: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=EMPTY; end
      16'd593: begin digit0<=THREE; digit1<=NINE; digit2<=FIVE; digit3<=EMPTY; end
      16'd594: begin digit0<=FOUR; digit1<=NINE; digit2<=FIVE; digit3<=EMPTY; end
      16'd595: begin digit0<=FIVE; digit1<=NINE; digit2<=FIVE; digit3<=EMPTY; end
      16'd596: begin digit0<=SIX; digit1<=NINE; digit2<=FIVE; digit3<=EMPTY; end
      16'd597: begin digit0<=SEVEN; digit1<=NINE; digit2<=FIVE; digit3<=EMPTY; end
      16'd598: begin digit0<=EIGHT; digit1<=NINE; digit2<=FIVE; digit3<=EMPTY; end
      16'd599: begin digit0<=NINE; digit1<=NINE; digit2<=FIVE; digit3<=EMPTY; end
	  16'd600: begin digit0<=ZERO; digit1<=ZERO; digit2<=SIX; digit3<=EMPTY; end
      16'd601: begin digit0<=ONE; digit1<=ZERO; digit2<=SIX; digit3<=EMPTY; end
      16'd602: begin digit0<=TWO; digit1<=ZERO; digit2<=SIX; digit3<=EMPTY; end
      16'd603: begin digit0<=THREE; digit1<=ZERO; digit2<=SIX; digit3<=EMPTY; end
      16'd604: begin digit0<=FOUR; digit1<=ZERO; digit2<=SIX; digit3<=EMPTY; end
      16'd605: begin digit0<=FIVE; digit1<=ZERO; digit2<=SIX; digit3<=EMPTY; end
      16'd606: begin digit0<=SIX; digit1<=ZERO; digit2<=SIX; digit3<=EMPTY; end
      16'd607: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SIX; digit3<=EMPTY; end
      16'd608: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SIX; digit3<=EMPTY; end
      16'd609: begin digit0<=NINE; digit1<=ZERO; digit2<=SIX; digit3<=EMPTY; end
      16'd610: begin digit0<=ZERO; digit1<=ONE; digit2<=SIX; digit3<=EMPTY; end
      16'd611: begin digit0<=ONE; digit1<=ONE; digit2<=SIX; digit3<=EMPTY; end
      16'd612: begin digit0<=TWO; digit1<=ONE; digit2<=SIX; digit3<=EMPTY; end
      16'd613: begin digit0<=THREE; digit1<=ONE; digit2<=SIX; digit3<=EMPTY; end
      16'd614: begin digit0<=FOUR; digit1<=ONE; digit2<=SIX; digit3<=EMPTY; end
      16'd615: begin digit0<=FIVE; digit1<=ONE; digit2<=SIX; digit3<=EMPTY; end
      16'd616: begin digit0<=SIX; digit1<=ONE; digit2<=SIX; digit3<=EMPTY; end
      16'd617: begin digit0<=SEVEN; digit1<=ONE; digit2<=SIX; digit3<=EMPTY; end
      16'd618: begin digit0<=EIGHT; digit1<=ONE; digit2<=SIX; digit3<=EMPTY; end
      16'd619: begin digit0<=NINE; digit1<=ONE; digit2<=SIX; digit3<=EMPTY; end
      16'd620: begin digit0<=ZERO; digit1<=TWO; digit2<=SIX; digit3<=EMPTY; end
      16'd621: begin digit0<=ONE; digit1<=TWO; digit2<=SIX; digit3<=EMPTY; end
      16'd622: begin digit0<=TWO; digit1<=TWO; digit2<=SIX; digit3<=EMPTY; end
      16'd623: begin digit0<=THREE; digit1<=TWO; digit2<=SIX; digit3<=EMPTY; end
      16'd624: begin digit0<=FOUR; digit1<=TWO; digit2<=SIX; digit3<=EMPTY; end
      16'd625: begin digit0<=FIVE; digit1<=TWO; digit2<=SIX; digit3<=EMPTY; end
      16'd626: begin digit0<=SIX; digit1<=TWO; digit2<=SIX; digit3<=EMPTY; end
      16'd627: begin digit0<=SEVEN; digit1<=TWO; digit2<=SIX; digit3<=EMPTY; end
      16'd628: begin digit0<=EIGHT; digit1<=TWO; digit2<=SIX; digit3<=EMPTY; end
      16'd629: begin digit0<=NINE; digit1<=TWO; digit2<=SIX; digit3<=EMPTY; end
      16'd630: begin digit0<=ZERO; digit1<=THREE; digit2<=SIX; digit3<=EMPTY; end
      16'd631: begin digit0<=ONE; digit1<=THREE; digit2<=SIX; digit3<=EMPTY; end
      16'd632: begin digit0<=TWO; digit1<=THREE; digit2<=SIX; digit3<=EMPTY; end
      16'd633: begin digit0<=THREE; digit1<=THREE; digit2<=SIX; digit3<=EMPTY; end
      16'd634: begin digit0<=FOUR; digit1<=THREE; digit2<=SIX; digit3<=EMPTY; end
      16'd635: begin digit0<=FIVE; digit1<=THREE; digit2<=SIX; digit3<=EMPTY; end
      16'd636: begin digit0<=SIX; digit1<=THREE; digit2<=SIX; digit3<=EMPTY; end
      16'd637: begin digit0<=SEVEN; digit1<=THREE; digit2<=SIX; digit3<=EMPTY; end
      16'd638: begin digit0<=EIGHT; digit1<=THREE; digit2<=SIX; digit3<=EMPTY; end
      16'd639: begin digit0<=NINE; digit1<=THREE; digit2<=SIX; digit3<=EMPTY; end
      16'd640: begin digit0<=ZERO; digit1<=FOUR; digit2<=SIX; digit3<=EMPTY; end
      16'd641: begin digit0<=ONE; digit1<=FOUR; digit2<=SIX; digit3<=EMPTY; end
      16'd642: begin digit0<=TWO; digit1<=FOUR; digit2<=SIX; digit3<=EMPTY; end
      16'd643: begin digit0<=THREE; digit1<=FOUR; digit2<=SIX; digit3<=EMPTY; end
      16'd644: begin digit0<=FOUR; digit1<=FOUR; digit2<=SIX; digit3<=EMPTY; end
      16'd645: begin digit0<=FIVE; digit1<=FOUR; digit2<=SIX; digit3<=EMPTY; end
      16'd646: begin digit0<=SIX; digit1<=FOUR; digit2<=SIX; digit3<=EMPTY; end
      16'd647: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SIX; digit3<=EMPTY; end
      16'd648: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SIX; digit3<=EMPTY; end
      16'd649: begin digit0<=NINE; digit1<=FOUR; digit2<=SIX; digit3<=EMPTY; end
      16'd650: begin digit0<=ZERO; digit1<=FIVE; digit2<=SIX; digit3<=EMPTY; end
      16'd651: begin digit0<=ONE; digit1<=FIVE; digit2<=SIX; digit3<=EMPTY; end
      16'd652: begin digit0<=TWO; digit1<=FIVE; digit2<=SIX; digit3<=EMPTY; end
      16'd653: begin digit0<=THREE; digit1<=FIVE; digit2<=SIX; digit3<=EMPTY; end
      16'd654: begin digit0<=FOUR; digit1<=FIVE; digit2<=SIX; digit3<=EMPTY; end
      16'd655: begin digit0<=FIVE; digit1<=FIVE; digit2<=SIX; digit3<=EMPTY; end
      16'd656: begin digit0<=SIX; digit1<=FIVE; digit2<=SIX; digit3<=EMPTY; end
      16'd657: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SIX; digit3<=EMPTY; end
      16'd658: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SIX; digit3<=EMPTY; end
      16'd659: begin digit0<=NINE; digit1<=FIVE; digit2<=SIX; digit3<=EMPTY; end
      16'd660: begin digit0<=ZERO; digit1<=SIX; digit2<=SIX; digit3<=EMPTY; end
      16'd661: begin digit0<=ONE; digit1<=SIX; digit2<=SIX; digit3<=EMPTY; end
      16'd662: begin digit0<=TWO; digit1<=SIX; digit2<=SIX; digit3<=EMPTY; end
      16'd663: begin digit0<=THREE; digit1<=SIX; digit2<=SIX; digit3<=EMPTY; end
      16'd664: begin digit0<=FOUR; digit1<=SIX; digit2<=SIX; digit3<=EMPTY; end
      16'd665: begin digit0<=FIVE; digit1<=SIX; digit2<=SIX; digit3<=EMPTY; end
      16'd666: begin digit0<=SIX; digit1<=SIX; digit2<=SIX; digit3<=EMPTY; end
      16'd667: begin digit0<=SEVEN; digit1<=SIX; digit2<=SIX; digit3<=EMPTY; end
      16'd668: begin digit0<=EIGHT; digit1<=SIX; digit2<=SIX; digit3<=EMPTY; end
      16'd669: begin digit0<=NINE; digit1<=SIX; digit2<=SIX; digit3<=EMPTY; end
      16'd670: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SIX; digit3<=EMPTY; end
      16'd671: begin digit0<=ONE; digit1<=SEVEN; digit2<=SIX; digit3<=EMPTY; end
      16'd672: begin digit0<=TWO; digit1<=SEVEN; digit2<=SIX; digit3<=EMPTY; end
      16'd673: begin digit0<=THREE; digit1<=SEVEN; digit2<=SIX; digit3<=EMPTY; end
      16'd674: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SIX; digit3<=EMPTY; end
      16'd675: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SIX; digit3<=EMPTY; end
      16'd676: begin digit0<=SIX; digit1<=SEVEN; digit2<=SIX; digit3<=EMPTY; end
      16'd677: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SIX; digit3<=EMPTY; end
      16'd678: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SIX; digit3<=EMPTY; end
      16'd679: begin digit0<=NINE; digit1<=SEVEN; digit2<=SIX; digit3<=EMPTY; end
      16'd680: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=EMPTY; end
      16'd681: begin digit0<=ONE; digit1<=EIGHT; digit2<=SIX; digit3<=EMPTY; end
      16'd682: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=EMPTY; end
      16'd683: begin digit0<=THREE; digit1<=EIGHT; digit2<=SIX; digit3<=EMPTY; end
      16'd684: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SIX; digit3<=EMPTY; end
      16'd685: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SIX; digit3<=EMPTY; end
      16'd686: begin digit0<=SIX; digit1<=EIGHT; digit2<=SIX; digit3<=EMPTY; end
      16'd687: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SIX; digit3<=EMPTY; end
      16'd688: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SIX; digit3<=EMPTY; end
      16'd689: begin digit0<=NINE; digit1<=EIGHT; digit2<=SIX; digit3<=EMPTY; end
      16'd690: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=EMPTY; end
      16'd691: begin digit0<=ONE; digit1<=NINE; digit2<=SIX; digit3<=EMPTY; end
      16'd692: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=EMPTY; end
      16'd693: begin digit0<=THREE; digit1<=NINE; digit2<=SIX; digit3<=EMPTY; end
      16'd694: begin digit0<=FOUR; digit1<=NINE; digit2<=SIX; digit3<=EMPTY; end
      16'd695: begin digit0<=FIVE; digit1<=NINE; digit2<=SIX; digit3<=EMPTY; end
      16'd696: begin digit0<=SIX; digit1<=NINE; digit2<=SIX; digit3<=EMPTY; end
      16'd697: begin digit0<=SEVEN; digit1<=NINE; digit2<=SIX; digit3<=EMPTY; end
      16'd698: begin digit0<=EIGHT; digit1<=NINE; digit2<=SIX; digit3<=EMPTY; end
      16'd699: begin digit0<=NINE; digit1<=NINE; digit2<=SIX; digit3<=EMPTY; end
	  16'd700: begin digit0<=ZERO; digit1<=ZERO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd701: begin digit0<=ONE; digit1<=ZERO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd702: begin digit0<=TWO; digit1<=ZERO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd703: begin digit0<=THREE; digit1<=ZERO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd704: begin digit0<=FOUR; digit1<=ZERO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd705: begin digit0<=FIVE; digit1<=ZERO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd706: begin digit0<=SIX; digit1<=ZERO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd707: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd708: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd709: begin digit0<=NINE; digit1<=ZERO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd710: begin digit0<=ZERO; digit1<=ONE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd711: begin digit0<=ONE; digit1<=ONE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd712: begin digit0<=TWO; digit1<=ONE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd713: begin digit0<=THREE; digit1<=ONE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd714: begin digit0<=FOUR; digit1<=ONE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd715: begin digit0<=FIVE; digit1<=ONE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd716: begin digit0<=SIX; digit1<=ONE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd717: begin digit0<=SEVEN; digit1<=ONE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd718: begin digit0<=EIGHT; digit1<=ONE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd719: begin digit0<=NINE; digit1<=ONE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd720: begin digit0<=ZERO; digit1<=TWO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd721: begin digit0<=ONE; digit1<=TWO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd722: begin digit0<=TWO; digit1<=TWO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd723: begin digit0<=THREE; digit1<=TWO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd724: begin digit0<=FOUR; digit1<=TWO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd725: begin digit0<=FIVE; digit1<=TWO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd726: begin digit0<=SIX; digit1<=TWO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd727: begin digit0<=SEVEN; digit1<=TWO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd728: begin digit0<=EIGHT; digit1<=TWO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd729: begin digit0<=NINE; digit1<=TWO; digit2<=SEVEN; digit3<=EMPTY; end
      16'd730: begin digit0<=ZERO; digit1<=THREE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd731: begin digit0<=ONE; digit1<=THREE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd732: begin digit0<=TWO; digit1<=THREE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd733: begin digit0<=THREE; digit1<=THREE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd734: begin digit0<=FOUR; digit1<=THREE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd735: begin digit0<=FIVE; digit1<=THREE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd736: begin digit0<=SIX; digit1<=THREE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd737: begin digit0<=SEVEN; digit1<=THREE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd738: begin digit0<=EIGHT; digit1<=THREE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd739: begin digit0<=NINE; digit1<=THREE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd740: begin digit0<=ZERO; digit1<=FOUR; digit2<=SEVEN; digit3<=EMPTY; end
      16'd741: begin digit0<=ONE; digit1<=FOUR; digit2<=SEVEN; digit3<=EMPTY; end
      16'd742: begin digit0<=TWO; digit1<=FOUR; digit2<=SEVEN; digit3<=EMPTY; end
      16'd743: begin digit0<=THREE; digit1<=FOUR; digit2<=SEVEN; digit3<=EMPTY; end
      16'd744: begin digit0<=FOUR; digit1<=FOUR; digit2<=SEVEN; digit3<=EMPTY; end
      16'd745: begin digit0<=FIVE; digit1<=FOUR; digit2<=SEVEN; digit3<=EMPTY; end
      16'd746: begin digit0<=SIX; digit1<=FOUR; digit2<=SEVEN; digit3<=EMPTY; end
      16'd747: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SEVEN; digit3<=EMPTY; end
      16'd748: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SEVEN; digit3<=EMPTY; end
      16'd749: begin digit0<=NINE; digit1<=FOUR; digit2<=SEVEN; digit3<=EMPTY; end
      16'd750: begin digit0<=ZERO; digit1<=FIVE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd751: begin digit0<=ONE; digit1<=FIVE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd752: begin digit0<=TWO; digit1<=FIVE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd753: begin digit0<=THREE; digit1<=FIVE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd754: begin digit0<=FOUR; digit1<=FIVE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd755: begin digit0<=FIVE; digit1<=FIVE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd756: begin digit0<=SIX; digit1<=FIVE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd757: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd758: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd759: begin digit0<=NINE; digit1<=FIVE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd760: begin digit0<=ZERO; digit1<=SIX; digit2<=SEVEN; digit3<=EMPTY; end
      16'd761: begin digit0<=ONE; digit1<=SIX; digit2<=SEVEN; digit3<=EMPTY; end
      16'd762: begin digit0<=TWO; digit1<=SIX; digit2<=SEVEN; digit3<=EMPTY; end
      16'd763: begin digit0<=THREE; digit1<=SIX; digit2<=SEVEN; digit3<=EMPTY; end
      16'd764: begin digit0<=FOUR; digit1<=SIX; digit2<=SEVEN; digit3<=EMPTY; end
      16'd765: begin digit0<=FIVE; digit1<=SIX; digit2<=SEVEN; digit3<=EMPTY; end
      16'd766: begin digit0<=SIX; digit1<=SIX; digit2<=SEVEN; digit3<=EMPTY; end
      16'd767: begin digit0<=SEVEN; digit1<=SIX; digit2<=SEVEN; digit3<=EMPTY; end
      16'd768: begin digit0<=EIGHT; digit1<=SIX; digit2<=SEVEN; digit3<=EMPTY; end
      16'd769: begin digit0<=NINE; digit1<=SIX; digit2<=SEVEN; digit3<=EMPTY; end
      16'd770: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SEVEN; digit3<=EMPTY; end
      16'd771: begin digit0<=ONE; digit1<=SEVEN; digit2<=SEVEN; digit3<=EMPTY; end
      16'd772: begin digit0<=TWO; digit1<=SEVEN; digit2<=SEVEN; digit3<=EMPTY; end
      16'd773: begin digit0<=THREE; digit1<=SEVEN; digit2<=SEVEN; digit3<=EMPTY; end
      16'd774: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SEVEN; digit3<=EMPTY; end
      16'd775: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SEVEN; digit3<=EMPTY; end
      16'd776: begin digit0<=SIX; digit1<=SEVEN; digit2<=SEVEN; digit3<=EMPTY; end
      16'd777: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SEVEN; digit3<=EMPTY; end
      16'd778: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SEVEN; digit3<=EMPTY; end
      16'd779: begin digit0<=NINE; digit1<=SEVEN; digit2<=SEVEN; digit3<=EMPTY; end
      16'd780: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=EMPTY; end
      16'd781: begin digit0<=ONE; digit1<=EIGHT; digit2<=SEVEN; digit3<=EMPTY; end
      16'd782: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=EMPTY; end
      16'd783: begin digit0<=THREE; digit1<=EIGHT; digit2<=SEVEN; digit3<=EMPTY; end
      16'd784: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SEVEN; digit3<=EMPTY; end
      16'd785: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SEVEN; digit3<=EMPTY; end
      16'd786: begin digit0<=SIX; digit1<=EIGHT; digit2<=SEVEN; digit3<=EMPTY; end
      16'd787: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SEVEN; digit3<=EMPTY; end
      16'd788: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SEVEN; digit3<=EMPTY; end
      16'd789: begin digit0<=NINE; digit1<=EIGHT; digit2<=SEVEN; digit3<=EMPTY; end
      16'd790: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd791: begin digit0<=ONE; digit1<=NINE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd792: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd793: begin digit0<=THREE; digit1<=NINE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd794: begin digit0<=FOUR; digit1<=NINE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd795: begin digit0<=FIVE; digit1<=NINE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd796: begin digit0<=SIX; digit1<=NINE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd797: begin digit0<=SEVEN; digit1<=NINE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd798: begin digit0<=EIGHT; digit1<=NINE; digit2<=SEVEN; digit3<=EMPTY; end
      16'd799: begin digit0<=NINE; digit1<=NINE; digit2<=SEVEN; digit3<=EMPTY; end
	  16'd800: begin digit0<=ZERO; digit1<=ZERO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd801: begin digit0<=ONE; digit1<=ZERO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd802: begin digit0<=TWO; digit1<=ZERO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd803: begin digit0<=THREE; digit1<=ZERO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd804: begin digit0<=FOUR; digit1<=ZERO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd805: begin digit0<=FIVE; digit1<=ZERO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd806: begin digit0<=SIX; digit1<=ZERO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd807: begin digit0<=SEVEN; digit1<=ZERO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd808: begin digit0<=EIGHT; digit1<=ZERO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd809: begin digit0<=NINE; digit1<=ZERO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd810: begin digit0<=ZERO; digit1<=ONE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd811: begin digit0<=ONE; digit1<=ONE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd812: begin digit0<=TWO; digit1<=ONE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd813: begin digit0<=THREE; digit1<=ONE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd814: begin digit0<=FOUR; digit1<=ONE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd815: begin digit0<=FIVE; digit1<=ONE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd816: begin digit0<=SIX; digit1<=ONE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd817: begin digit0<=SEVEN; digit1<=ONE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd818: begin digit0<=EIGHT; digit1<=ONE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd819: begin digit0<=NINE; digit1<=ONE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd820: begin digit0<=ZERO; digit1<=TWO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd821: begin digit0<=ONE; digit1<=TWO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd822: begin digit0<=TWO; digit1<=TWO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd823: begin digit0<=THREE; digit1<=TWO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd824: begin digit0<=FOUR; digit1<=TWO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd825: begin digit0<=FIVE; digit1<=TWO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd826: begin digit0<=SIX; digit1<=TWO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd827: begin digit0<=SEVEN; digit1<=TWO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd828: begin digit0<=EIGHT; digit1<=TWO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd829: begin digit0<=NINE; digit1<=TWO; digit2<=EIGHT; digit3<=EMPTY; end
      16'd830: begin digit0<=ZERO; digit1<=THREE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd831: begin digit0<=ONE; digit1<=THREE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd832: begin digit0<=TWO; digit1<=THREE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd833: begin digit0<=THREE; digit1<=THREE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd834: begin digit0<=FOUR; digit1<=THREE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd835: begin digit0<=FIVE; digit1<=THREE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd836: begin digit0<=SIX; digit1<=THREE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd837: begin digit0<=SEVEN; digit1<=THREE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd838: begin digit0<=EIGHT; digit1<=THREE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd839: begin digit0<=NINE; digit1<=THREE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd840: begin digit0<=ZERO; digit1<=FOUR; digit2<=EIGHT; digit3<=EMPTY; end
      16'd841: begin digit0<=ONE; digit1<=FOUR; digit2<=EIGHT; digit3<=EMPTY; end
      16'd842: begin digit0<=TWO; digit1<=FOUR; digit2<=EIGHT; digit3<=EMPTY; end
      16'd843: begin digit0<=THREE; digit1<=FOUR; digit2<=EIGHT; digit3<=EMPTY; end
      16'd844: begin digit0<=FOUR; digit1<=FOUR; digit2<=EIGHT; digit3<=EMPTY; end
      16'd845: begin digit0<=FIVE; digit1<=FOUR; digit2<=EIGHT; digit3<=EMPTY; end
      16'd846: begin digit0<=SIX; digit1<=FOUR; digit2<=EIGHT; digit3<=EMPTY; end
      16'd847: begin digit0<=SEVEN; digit1<=FOUR; digit2<=EIGHT; digit3<=EMPTY; end
      16'd848: begin digit0<=EIGHT; digit1<=FOUR; digit2<=EIGHT; digit3<=EMPTY; end
      16'd849: begin digit0<=NINE; digit1<=FOUR; digit2<=EIGHT; digit3<=EMPTY; end
      16'd850: begin digit0<=ZERO; digit1<=FIVE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd851: begin digit0<=ONE; digit1<=FIVE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd852: begin digit0<=TWO; digit1<=FIVE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd853: begin digit0<=THREE; digit1<=FIVE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd854: begin digit0<=FOUR; digit1<=FIVE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd855: begin digit0<=FIVE; digit1<=FIVE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd856: begin digit0<=SIX; digit1<=FIVE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd857: begin digit0<=SEVEN; digit1<=FIVE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd858: begin digit0<=EIGHT; digit1<=FIVE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd859: begin digit0<=NINE; digit1<=FIVE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd860: begin digit0<=ZERO; digit1<=SIX; digit2<=EIGHT; digit3<=EMPTY; end
      16'd861: begin digit0<=ONE; digit1<=SIX; digit2<=EIGHT; digit3<=EMPTY; end
      16'd862: begin digit0<=TWO; digit1<=SIX; digit2<=EIGHT; digit3<=EMPTY; end
      16'd863: begin digit0<=THREE; digit1<=SIX; digit2<=EIGHT; digit3<=EMPTY; end
      16'd864: begin digit0<=FOUR; digit1<=SIX; digit2<=EIGHT; digit3<=EMPTY; end
      16'd865: begin digit0<=FIVE; digit1<=SIX; digit2<=EIGHT; digit3<=EMPTY; end
      16'd866: begin digit0<=SIX; digit1<=SIX; digit2<=EIGHT; digit3<=EMPTY; end
      16'd867: begin digit0<=SEVEN; digit1<=SIX; digit2<=EIGHT; digit3<=EMPTY; end
      16'd868: begin digit0<=EIGHT; digit1<=SIX; digit2<=EIGHT; digit3<=EMPTY; end
      16'd869: begin digit0<=NINE; digit1<=SIX; digit2<=EIGHT; digit3<=EMPTY; end
      16'd870: begin digit0<=ZERO; digit1<=SEVEN; digit2<=EIGHT; digit3<=EMPTY; end
      16'd871: begin digit0<=ONE; digit1<=SEVEN; digit2<=EIGHT; digit3<=EMPTY; end
      16'd872: begin digit0<=TWO; digit1<=SEVEN; digit2<=EIGHT; digit3<=EMPTY; end
      16'd873: begin digit0<=THREE; digit1<=SEVEN; digit2<=EIGHT; digit3<=EMPTY; end
      16'd874: begin digit0<=FOUR; digit1<=SEVEN; digit2<=EIGHT; digit3<=EMPTY; end
      16'd875: begin digit0<=FIVE; digit1<=SEVEN; digit2<=EIGHT; digit3<=EMPTY; end
      16'd876: begin digit0<=SIX; digit1<=SEVEN; digit2<=EIGHT; digit3<=EMPTY; end
      16'd877: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=EIGHT; digit3<=EMPTY; end
      16'd878: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=EIGHT; digit3<=EMPTY; end
      16'd879: begin digit0<=NINE; digit1<=SEVEN; digit2<=EIGHT; digit3<=EMPTY; end
      16'd880: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=EMPTY; end
      16'd881: begin digit0<=ONE; digit1<=EIGHT; digit2<=EIGHT; digit3<=EMPTY; end
      16'd882: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=EMPTY; end
      16'd883: begin digit0<=THREE; digit1<=EIGHT; digit2<=EIGHT; digit3<=EMPTY; end
      16'd884: begin digit0<=FOUR; digit1<=EIGHT; digit2<=EIGHT; digit3<=EMPTY; end
      16'd885: begin digit0<=FIVE; digit1<=EIGHT; digit2<=EIGHT; digit3<=EMPTY; end
      16'd886: begin digit0<=SIX; digit1<=EIGHT; digit2<=EIGHT; digit3<=EMPTY; end
      16'd887: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=EIGHT; digit3<=EMPTY; end
      16'd888: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=EIGHT; digit3<=EMPTY; end
      16'd889: begin digit0<=NINE; digit1<=EIGHT; digit2<=EIGHT; digit3<=EMPTY; end
      16'd890: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd891: begin digit0<=ONE; digit1<=NINE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd892: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd893: begin digit0<=THREE; digit1<=NINE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd894: begin digit0<=FOUR; digit1<=NINE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd895: begin digit0<=FIVE; digit1<=NINE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd896: begin digit0<=SIX; digit1<=NINE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd897: begin digit0<=SEVEN; digit1<=NINE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd898: begin digit0<=EIGHT; digit1<=NINE; digit2<=EIGHT; digit3<=EMPTY; end
      16'd899: begin digit0<=NINE; digit1<=NINE; digit2<=EIGHT; digit3<=EMPTY; end
	  16'd900: begin digit0<=ZERO; digit1<=ZERO; digit2<=NINE; digit3<=EMPTY; end
      16'd901: begin digit0<=ONE; digit1<=ZERO; digit2<=NINE; digit3<=EMPTY; end
      16'd902: begin digit0<=TWO; digit1<=ZERO; digit2<=NINE; digit3<=EMPTY; end
      16'd903: begin digit0<=THREE; digit1<=ZERO; digit2<=NINE; digit3<=EMPTY; end
      16'd904: begin digit0<=FOUR; digit1<=ZERO; digit2<=NINE; digit3<=EMPTY; end
      16'd905: begin digit0<=FIVE; digit1<=ZERO; digit2<=NINE; digit3<=EMPTY; end
      16'd906: begin digit0<=SIX; digit1<=ZERO; digit2<=NINE; digit3<=EMPTY; end
      16'd907: begin digit0<=SEVEN; digit1<=ZERO; digit2<=NINE; digit3<=EMPTY; end
      16'd908: begin digit0<=EIGHT; digit1<=ZERO; digit2<=NINE; digit3<=EMPTY; end
      16'd909: begin digit0<=NINE; digit1<=ZERO; digit2<=NINE; digit3<=EMPTY; end
      16'd910: begin digit0<=ZERO; digit1<=ONE; digit2<=NINE; digit3<=EMPTY; end
      16'd911: begin digit0<=ONE; digit1<=ONE; digit2<=NINE; digit3<=EMPTY; end
      16'd912: begin digit0<=TWO; digit1<=ONE; digit2<=NINE; digit3<=EMPTY; end
      16'd913: begin digit0<=THREE; digit1<=ONE; digit2<=NINE; digit3<=EMPTY; end
      16'd914: begin digit0<=FOUR; digit1<=ONE; digit2<=NINE; digit3<=EMPTY; end
      16'd915: begin digit0<=FIVE; digit1<=ONE; digit2<=NINE; digit3<=EMPTY; end
      16'd916: begin digit0<=SIX; digit1<=ONE; digit2<=NINE; digit3<=EMPTY; end
      16'd917: begin digit0<=SEVEN; digit1<=ONE; digit2<=NINE; digit3<=EMPTY; end
      16'd918: begin digit0<=EIGHT; digit1<=ONE; digit2<=NINE; digit3<=EMPTY; end
      16'd919: begin digit0<=NINE; digit1<=ONE; digit2<=NINE; digit3<=EMPTY; end
      16'd920: begin digit0<=ZERO; digit1<=TWO; digit2<=NINE; digit3<=EMPTY; end
      16'd921: begin digit0<=ONE; digit1<=TWO; digit2<=NINE; digit3<=EMPTY; end
      16'd922: begin digit0<=TWO; digit1<=TWO; digit2<=NINE; digit3<=EMPTY; end
      16'd923: begin digit0<=THREE; digit1<=TWO; digit2<=NINE; digit3<=EMPTY; end
      16'd924: begin digit0<=FOUR; digit1<=TWO; digit2<=NINE; digit3<=EMPTY; end
      16'd925: begin digit0<=FIVE; digit1<=TWO; digit2<=NINE; digit3<=EMPTY; end
      16'd926: begin digit0<=SIX; digit1<=TWO; digit2<=NINE; digit3<=EMPTY; end
      16'd927: begin digit0<=SEVEN; digit1<=TWO; digit2<=NINE; digit3<=EMPTY; end
      16'd928: begin digit0<=EIGHT; digit1<=TWO; digit2<=NINE; digit3<=EMPTY; end
      16'd929: begin digit0<=NINE; digit1<=TWO; digit2<=NINE; digit3<=EMPTY; end
      16'd930: begin digit0<=ZERO; digit1<=THREE; digit2<=NINE; digit3<=EMPTY; end
      16'd931: begin digit0<=ONE; digit1<=THREE; digit2<=NINE; digit3<=EMPTY; end
      16'd932: begin digit0<=TWO; digit1<=THREE; digit2<=NINE; digit3<=EMPTY; end
      16'd933: begin digit0<=THREE; digit1<=THREE; digit2<=NINE; digit3<=EMPTY; end
      16'd934: begin digit0<=FOUR; digit1<=THREE; digit2<=NINE; digit3<=EMPTY; end
      16'd935: begin digit0<=FIVE; digit1<=THREE; digit2<=NINE; digit3<=EMPTY; end
      16'd936: begin digit0<=SIX; digit1<=THREE; digit2<=NINE; digit3<=EMPTY; end
      16'd937: begin digit0<=SEVEN; digit1<=THREE; digit2<=NINE; digit3<=EMPTY; end
      16'd938: begin digit0<=EIGHT; digit1<=THREE; digit2<=NINE; digit3<=EMPTY; end
      16'd939: begin digit0<=NINE; digit1<=THREE; digit2<=NINE; digit3<=EMPTY; end
      16'd940: begin digit0<=ZERO; digit1<=FOUR; digit2<=NINE; digit3<=EMPTY; end
      16'd941: begin digit0<=ONE; digit1<=FOUR; digit2<=NINE; digit3<=EMPTY; end
      16'd942: begin digit0<=TWO; digit1<=FOUR; digit2<=NINE; digit3<=EMPTY; end
      16'd943: begin digit0<=THREE; digit1<=FOUR; digit2<=NINE; digit3<=EMPTY; end
      16'd944: begin digit0<=FOUR; digit1<=FOUR; digit2<=NINE; digit3<=EMPTY; end
      16'd945: begin digit0<=FIVE; digit1<=FOUR; digit2<=NINE; digit3<=EMPTY; end
      16'd946: begin digit0<=SIX; digit1<=FOUR; digit2<=NINE; digit3<=EMPTY; end
      16'd947: begin digit0<=SEVEN; digit1<=FOUR; digit2<=NINE; digit3<=EMPTY; end
      16'd948: begin digit0<=EIGHT; digit1<=FOUR; digit2<=NINE; digit3<=EMPTY; end
      16'd949: begin digit0<=NINE; digit1<=FOUR; digit2<=NINE; digit3<=EMPTY; end
      16'd950: begin digit0<=ZERO; digit1<=FIVE; digit2<=NINE; digit3<=EMPTY; end
      16'd951: begin digit0<=ONE; digit1<=FIVE; digit2<=NINE; digit3<=EMPTY; end
      16'd952: begin digit0<=TWO; digit1<=FIVE; digit2<=NINE; digit3<=EMPTY; end
      16'd953: begin digit0<=THREE; digit1<=FIVE; digit2<=NINE; digit3<=EMPTY; end
      16'd954: begin digit0<=FOUR; digit1<=FIVE; digit2<=NINE; digit3<=EMPTY; end
      16'd955: begin digit0<=FIVE; digit1<=FIVE; digit2<=NINE; digit3<=EMPTY; end
      16'd956: begin digit0<=SIX; digit1<=FIVE; digit2<=NINE; digit3<=EMPTY; end
      16'd957: begin digit0<=SEVEN; digit1<=FIVE; digit2<=NINE; digit3<=EMPTY; end
      16'd958: begin digit0<=EIGHT; digit1<=FIVE; digit2<=NINE; digit3<=EMPTY; end
      16'd959: begin digit0<=NINE; digit1<=FIVE; digit2<=NINE; digit3<=EMPTY; end
      16'd960: begin digit0<=ZERO; digit1<=SIX; digit2<=NINE; digit3<=EMPTY; end
      16'd961: begin digit0<=ONE; digit1<=SIX; digit2<=NINE; digit3<=EMPTY; end
      16'd962: begin digit0<=TWO; digit1<=SIX; digit2<=NINE; digit3<=EMPTY; end
      16'd963: begin digit0<=THREE; digit1<=SIX; digit2<=NINE; digit3<=EMPTY; end
      16'd964: begin digit0<=FOUR; digit1<=SIX; digit2<=NINE; digit3<=EMPTY; end
      16'd965: begin digit0<=FIVE; digit1<=SIX; digit2<=NINE; digit3<=EMPTY; end
      16'd966: begin digit0<=SIX; digit1<=SIX; digit2<=NINE; digit3<=EMPTY; end
      16'd967: begin digit0<=SEVEN; digit1<=SIX; digit2<=NINE; digit3<=EMPTY; end
      16'd968: begin digit0<=EIGHT; digit1<=SIX; digit2<=NINE; digit3<=EMPTY; end
      16'd969: begin digit0<=NINE; digit1<=SIX; digit2<=NINE; digit3<=EMPTY; end
      16'd970: begin digit0<=ZERO; digit1<=SEVEN; digit2<=NINE; digit3<=EMPTY; end
      16'd971: begin digit0<=ONE; digit1<=SEVEN; digit2<=NINE; digit3<=EMPTY; end
      16'd972: begin digit0<=TWO; digit1<=SEVEN; digit2<=NINE; digit3<=EMPTY; end
      16'd973: begin digit0<=THREE; digit1<=SEVEN; digit2<=NINE; digit3<=EMPTY; end
      16'd974: begin digit0<=FOUR; digit1<=SEVEN; digit2<=NINE; digit3<=EMPTY; end
      16'd975: begin digit0<=FIVE; digit1<=SEVEN; digit2<=NINE; digit3<=EMPTY; end
      16'd976: begin digit0<=SIX; digit1<=SEVEN; digit2<=NINE; digit3<=EMPTY; end
      16'd977: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=NINE; digit3<=EMPTY; end
      16'd978: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=NINE; digit3<=EMPTY; end
      16'd979: begin digit0<=NINE; digit1<=SEVEN; digit2<=NINE; digit3<=EMPTY; end
      16'd980: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=EMPTY; end
      16'd981: begin digit0<=ONE; digit1<=EIGHT; digit2<=NINE; digit3<=EMPTY; end
      16'd982: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=EMPTY; end
      16'd983: begin digit0<=THREE; digit1<=EIGHT; digit2<=NINE; digit3<=EMPTY; end
      16'd984: begin digit0<=FOUR; digit1<=EIGHT; digit2<=NINE; digit3<=EMPTY; end
      16'd985: begin digit0<=FIVE; digit1<=EIGHT; digit2<=NINE; digit3<=EMPTY; end
      16'd986: begin digit0<=SIX; digit1<=EIGHT; digit2<=NINE; digit3<=EMPTY; end
      16'd987: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=NINE; digit3<=EMPTY; end
      16'd988: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=NINE; digit3<=EMPTY; end
      16'd989: begin digit0<=NINE; digit1<=EIGHT; digit2<=NINE; digit3<=EMPTY; end
      16'd990: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=EMPTY; end
      16'd991: begin digit0<=ONE; digit1<=NINE; digit2<=NINE; digit3<=EMPTY; end
      16'd992: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=EMPTY; end
      16'd993: begin digit0<=THREE; digit1<=NINE; digit2<=NINE; digit3<=EMPTY; end
      16'd994: begin digit0<=FOUR; digit1<=NINE; digit2<=NINE; digit3<=EMPTY; end
      16'd995: begin digit0<=FIVE; digit1<=NINE; digit2<=NINE; digit3<=EMPTY; end
      16'd996: begin digit0<=SIX; digit1<=NINE; digit2<=NINE; digit3<=EMPTY; end
      16'd997: begin digit0<=SEVEN; digit1<=NINE; digit2<=NINE; digit3<=EMPTY; end
      16'd998: begin digit0<=EIGHT; digit1<=NINE; digit2<=NINE; digit3<=EMPTY; end
      16'd999: begin digit0<=NINE; digit1<=NINE; digit2<=NINE; digit3<=EMPTY; end
	  16'd1000: begin digit0<=ZERO; digit1<=ZERO; digit2<=ZERO; digit3<=ONE; end
      16'd1001: begin digit0<=ONE; digit1<=ZERO; digit2<=ZERO; digit3<=ONE; end
      16'd1002: begin digit0<=TWO; digit1<=ZERO; digit2<=ZERO; digit3<=ONE; end
      16'd1003: begin digit0<=THREE; digit1<=ZERO; digit2<=ZERO; digit3<=ONE; end
      16'd1004: begin digit0<=FOUR; digit1<=ZERO; digit2<=ZERO; digit3<=ONE; end
      16'd1005: begin digit0<=FIVE; digit1<=ZERO; digit2<=ZERO; digit3<=ONE; end
      16'd1006: begin digit0<=SIX; digit1<=ZERO; digit2<=ZERO; digit3<=ONE; end
      16'd1007: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ZERO; digit3<=ONE; end
      16'd1008: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ZERO; digit3<=ONE; end
      16'd1009: begin digit0<=NINE; digit1<=ZERO; digit2<=ZERO; digit3<=ONE; end
      16'd1010: begin digit0<=ZERO; digit1<=ONE; digit2<=ZERO; digit3<=ONE; end
      16'd1011: begin digit0<=ONE; digit1<=ONE; digit2<=ZERO; digit3<=ONE; end
      16'd1012: begin digit0<=TWO; digit1<=ONE; digit2<=ZERO; digit3<=ONE; end
      16'd1013: begin digit0<=THREE; digit1<=ONE; digit2<=ZERO; digit3<=ONE; end
      16'd1014: begin digit0<=FOUR; digit1<=ONE; digit2<=ZERO; digit3<=ONE; end
      16'd1015: begin digit0<=FIVE; digit1<=ONE; digit2<=ZERO; digit3<=ONE; end
      16'd1016: begin digit0<=SIX; digit1<=ONE; digit2<=ZERO; digit3<=ONE; end
      16'd1017: begin digit0<=SEVEN; digit1<=ONE; digit2<=ZERO; digit3<=ONE; end
      16'd1018: begin digit0<=EIGHT; digit1<=ONE; digit2<=ZERO; digit3<=ONE; end
      16'd1019: begin digit0<=NINE; digit1<=ONE; digit2<=ZERO; digit3<=ONE; end
      16'd1020: begin digit0<=ZERO; digit1<=TWO; digit2<=ZERO; digit3<=ONE; end
      16'd1021: begin digit0<=ONE; digit1<=TWO; digit2<=ZERO; digit3<=ONE; end
      16'd1022: begin digit0<=TWO; digit1<=TWO; digit2<=ZERO; digit3<=ONE; end
      16'd1023: begin digit0<=THREE; digit1<=TWO; digit2<=ZERO; digit3<=ONE; end
      16'd1024: begin digit0<=FOUR; digit1<=TWO; digit2<=ZERO; digit3<=ONE; end
      16'd1025: begin digit0<=FIVE; digit1<=TWO; digit2<=ZERO; digit3<=ONE; end
      16'd1026: begin digit0<=SIX; digit1<=TWO; digit2<=ZERO; digit3<=ONE; end
      16'd1027: begin digit0<=SEVEN; digit1<=TWO; digit2<=ZERO; digit3<=ONE; end
      16'd1028: begin digit0<=EIGHT; digit1<=TWO; digit2<=ZERO; digit3<=ONE; end
      16'd1029: begin digit0<=NINE; digit1<=TWO; digit2<=ZERO; digit3<=ONE; end
      16'd1030: begin digit0<=ZERO; digit1<=THREE; digit2<=ZERO; digit3<=ONE; end
      16'd1031: begin digit0<=ONE; digit1<=THREE; digit2<=ZERO; digit3<=ONE; end
      16'd1032: begin digit0<=TWO; digit1<=THREE; digit2<=ZERO; digit3<=ONE; end
      16'd1033: begin digit0<=THREE; digit1<=THREE; digit2<=ZERO; digit3<=ONE; end
      16'd1034: begin digit0<=FOUR; digit1<=THREE; digit2<=ZERO; digit3<=ONE; end
      16'd1035: begin digit0<=FIVE; digit1<=THREE; digit2<=ZERO; digit3<=ONE; end
      16'd1036: begin digit0<=SIX; digit1<=THREE; digit2<=ZERO; digit3<=ONE; end
      16'd1037: begin digit0<=SEVEN; digit1<=THREE; digit2<=ZERO; digit3<=ONE; end
      16'd1038: begin digit0<=EIGHT; digit1<=THREE; digit2<=ZERO; digit3<=ONE; end
      16'd1039: begin digit0<=NINE; digit1<=THREE; digit2<=ZERO; digit3<=ONE; end
      16'd1040: begin digit0<=ZERO; digit1<=FOUR; digit2<=ZERO; digit3<=ONE; end
      16'd1041: begin digit0<=ONE; digit1<=FOUR; digit2<=ZERO; digit3<=ONE; end
      16'd1042: begin digit0<=TWO; digit1<=FOUR; digit2<=ZERO; digit3<=ONE; end
      16'd1043: begin digit0<=THREE; digit1<=FOUR; digit2<=ZERO; digit3<=ONE; end
      16'd1044: begin digit0<=FOUR; digit1<=FOUR; digit2<=ZERO; digit3<=ONE; end
      16'd1045: begin digit0<=FIVE; digit1<=FOUR; digit2<=ZERO; digit3<=ONE; end
      16'd1046: begin digit0<=SIX; digit1<=FOUR; digit2<=ZERO; digit3<=ONE; end
      16'd1047: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ZERO; digit3<=ONE; end
      16'd1048: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ZERO; digit3<=ONE; end
      16'd1049: begin digit0<=NINE; digit1<=FOUR; digit2<=ZERO; digit3<=ONE; end
      16'd1050: begin digit0<=ZERO; digit1<=FIVE; digit2<=ZERO; digit3<=ONE; end
      16'd1051: begin digit0<=ONE; digit1<=FIVE; digit2<=ZERO; digit3<=ONE; end
      16'd1052: begin digit0<=TWO; digit1<=FIVE; digit2<=ZERO; digit3<=ONE; end
      16'd1053: begin digit0<=THREE; digit1<=FIVE; digit2<=ZERO; digit3<=ONE; end
      16'd1054: begin digit0<=FOUR; digit1<=FIVE; digit2<=ZERO; digit3<=ONE; end
      16'd1055: begin digit0<=FIVE; digit1<=FIVE; digit2<=ZERO; digit3<=ONE; end
      16'd1056: begin digit0<=SIX; digit1<=FIVE; digit2<=ZERO; digit3<=ONE; end
      16'd1057: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ZERO; digit3<=ONE; end
      16'd1058: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ZERO; digit3<=ONE; end
      16'd1059: begin digit0<=NINE; digit1<=FIVE; digit2<=ZERO; digit3<=ONE; end
      16'd1060: begin digit0<=ZERO; digit1<=SIX; digit2<=ZERO; digit3<=ONE; end
      16'd1061: begin digit0<=ONE; digit1<=SIX; digit2<=ZERO; digit3<=ONE; end
      16'd1062: begin digit0<=TWO; digit1<=SIX; digit2<=ZERO; digit3<=ONE; end
      16'd1063: begin digit0<=THREE; digit1<=SIX; digit2<=ZERO; digit3<=ONE; end
      16'd1064: begin digit0<=FOUR; digit1<=SIX; digit2<=ZERO; digit3<=ONE; end
      16'd1065: begin digit0<=FIVE; digit1<=SIX; digit2<=ZERO; digit3<=ONE; end
      16'd1066: begin digit0<=SIX; digit1<=SIX; digit2<=ZERO; digit3<=ONE; end
      16'd1067: begin digit0<=SEVEN; digit1<=SIX; digit2<=ZERO; digit3<=ONE; end
      16'd1068: begin digit0<=EIGHT; digit1<=SIX; digit2<=ZERO; digit3<=ONE; end
      16'd1069: begin digit0<=NINE; digit1<=SIX; digit2<=ZERO; digit3<=ONE; end
      16'd1070: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ZERO; digit3<=ONE; end
      16'd1071: begin digit0<=ONE; digit1<=SEVEN; digit2<=ZERO; digit3<=ONE; end
      16'd1072: begin digit0<=TWO; digit1<=SEVEN; digit2<=ZERO; digit3<=ONE; end
      16'd1073: begin digit0<=THREE; digit1<=SEVEN; digit2<=ZERO; digit3<=ONE; end
      16'd1074: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ZERO; digit3<=ONE; end
      16'd1075: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ZERO; digit3<=ONE; end
      16'd1076: begin digit0<=SIX; digit1<=SEVEN; digit2<=ZERO; digit3<=ONE; end
      16'd1077: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ZERO; digit3<=ONE; end
      16'd1078: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ZERO; digit3<=ONE; end
      16'd1079: begin digit0<=NINE; digit1<=SEVEN; digit2<=ZERO; digit3<=ONE; end
      16'd1080: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ZERO; digit3<=ONE; end
      16'd1081: begin digit0<=ONE; digit1<=EIGHT; digit2<=ZERO; digit3<=ONE; end
      16'd1082: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ZERO; digit3<=ONE; end
      16'd1083: begin digit0<=THREE; digit1<=EIGHT; digit2<=ZERO; digit3<=ONE; end
      16'd1084: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ZERO; digit3<=ONE; end
      16'd1085: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ZERO; digit3<=ONE; end
      16'd1086: begin digit0<=SIX; digit1<=EIGHT; digit2<=ZERO; digit3<=ONE; end
      16'd1087: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ZERO; digit3<=ONE; end
      16'd1088: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ZERO; digit3<=ONE; end
      16'd1089: begin digit0<=NINE; digit1<=EIGHT; digit2<=ZERO; digit3<=ONE; end
      16'd1090: begin digit0<=ZERO; digit1<=NINE; digit2<=ZERO; digit3<=ONE; end
      16'd1091: begin digit0<=ONE; digit1<=NINE; digit2<=ZERO; digit3<=ONE; end
      16'd1092: begin digit0<=ZERO; digit1<=NINE; digit2<=ZERO; digit3<=ONE; end
      16'd1093: begin digit0<=THREE; digit1<=NINE; digit2<=ZERO; digit3<=ONE; end
      16'd1094: begin digit0<=FOUR; digit1<=NINE; digit2<=ZERO; digit3<=ONE; end
      16'd1095: begin digit0<=FIVE; digit1<=NINE; digit2<=ZERO; digit3<=ONE; end
      16'd1096: begin digit0<=SIX; digit1<=NINE; digit2<=ZERO; digit3<=ONE; end
      16'd1097: begin digit0<=SEVEN; digit1<=NINE; digit2<=ZERO; digit3<=ONE; end
      16'd1098: begin digit0<=EIGHT; digit1<=NINE; digit2<=ZERO; digit3<=ONE; end
      16'd1099: begin digit0<=NINE; digit1<=NINE; digit2<=ZERO; digit3<=ONE; end
	  16'd1100: begin digit0<=ZERO; digit1<=ZERO; digit2<=ONE; digit3<=ONE; end
      16'd1101: begin digit0<=ONE; digit1<=ZERO; digit2<=ONE; digit3<=ONE; end
      16'd1102: begin digit0<=TWO; digit1<=ZERO; digit2<=ONE; digit3<=ONE; end
      16'd1103: begin digit0<=THREE; digit1<=ZERO; digit2<=ONE; digit3<=ONE; end
      16'd1104: begin digit0<=FOUR; digit1<=ZERO; digit2<=ONE; digit3<=ONE; end
      16'd1105: begin digit0<=FIVE; digit1<=ZERO; digit2<=ONE; digit3<=ONE; end
      16'd1106: begin digit0<=SIX; digit1<=ZERO; digit2<=ONE; digit3<=ONE; end
      16'd1107: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ONE; digit3<=ONE; end
      16'd1108: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ONE; digit3<=ONE; end
      16'd1109: begin digit0<=NINE; digit1<=ZERO; digit2<=ONE; digit3<=ONE; end
      16'd1110: begin digit0<=ZERO; digit1<=ONE; digit2<=ONE; digit3<=ONE; end
      16'd1111: begin digit0<=ONE; digit1<=ONE; digit2<=ONE; digit3<=ONE; end
      16'd1112: begin digit0<=TWO; digit1<=ONE; digit2<=ONE; digit3<=ONE; end
      16'd1113: begin digit0<=THREE; digit1<=ONE; digit2<=ONE; digit3<=ONE; end
      16'd1114: begin digit0<=FOUR; digit1<=ONE; digit2<=ONE; digit3<=ONE; end
      16'd1115: begin digit0<=FIVE; digit1<=ONE; digit2<=ONE; digit3<=ONE; end
      16'd1116: begin digit0<=SIX; digit1<=ONE; digit2<=ONE; digit3<=ONE; end
      16'd1117: begin digit0<=SEVEN; digit1<=ONE; digit2<=ONE; digit3<=ONE; end
      16'd1118: begin digit0<=EIGHT; digit1<=ONE; digit2<=ONE; digit3<=ONE; end
      16'd1119: begin digit0<=NINE; digit1<=ONE; digit2<=ONE; digit3<=ONE; end
      16'd1120: begin digit0<=ZERO; digit1<=TWO; digit2<=ONE; digit3<=ONE; end
      16'd1121: begin digit0<=ONE; digit1<=TWO; digit2<=ONE; digit3<=ONE; end
      16'd1122: begin digit0<=TWO; digit1<=TWO; digit2<=ONE; digit3<=ONE; end
      16'd1123: begin digit0<=THREE; digit1<=TWO; digit2<=ONE; digit3<=ONE; end
      16'd1124: begin digit0<=FOUR; digit1<=TWO; digit2<=ONE; digit3<=ONE; end
      16'd1125: begin digit0<=FIVE; digit1<=TWO; digit2<=ONE; digit3<=ONE; end
      16'd1126: begin digit0<=SIX; digit1<=TWO; digit2<=ONE; digit3<=ONE; end
      16'd1127: begin digit0<=SEVEN; digit1<=TWO; digit2<=ONE; digit3<=ONE; end
      16'd1128: begin digit0<=EIGHT; digit1<=TWO; digit2<=ONE; digit3<=ONE; end
      16'd1129: begin digit0<=NINE; digit1<=TWO; digit2<=ONE; digit3<=ONE; end
      16'd1130: begin digit0<=ZERO; digit1<=THREE; digit2<=ONE; digit3<=ONE; end
      16'd1131: begin digit0<=ONE; digit1<=THREE; digit2<=ONE; digit3<=ONE; end
      16'd1132: begin digit0<=TWO; digit1<=THREE; digit2<=ONE; digit3<=ONE; end
      16'd1133: begin digit0<=THREE; digit1<=THREE; digit2<=ONE; digit3<=ONE; end
      16'd1134: begin digit0<=FOUR; digit1<=THREE; digit2<=ONE; digit3<=ONE; end
      16'd1135: begin digit0<=FIVE; digit1<=THREE; digit2<=ONE; digit3<=ONE; end
      16'd1136: begin digit0<=SIX; digit1<=THREE; digit2<=ONE; digit3<=ONE; end
      16'd1137: begin digit0<=SEVEN; digit1<=THREE; digit2<=ONE; digit3<=ONE; end
      16'd1138: begin digit0<=EIGHT; digit1<=THREE; digit2<=ONE; digit3<=ONE; end
      16'd1139: begin digit0<=NINE; digit1<=THREE; digit2<=ONE; digit3<=ONE; end
      16'd1140: begin digit0<=ZERO; digit1<=FOUR; digit2<=ONE; digit3<=ONE; end
      16'd1141: begin digit0<=ONE; digit1<=FOUR; digit2<=ONE; digit3<=ONE; end
      16'd1142: begin digit0<=TWO; digit1<=FOUR; digit2<=ONE; digit3<=ONE; end
      16'd1143: begin digit0<=THREE; digit1<=FOUR; digit2<=ONE; digit3<=ONE; end
      16'd1144: begin digit0<=FOUR; digit1<=FOUR; digit2<=ONE; digit3<=ONE; end
      16'd1145: begin digit0<=FIVE; digit1<=FOUR; digit2<=ONE; digit3<=ONE; end
      16'd1146: begin digit0<=SIX; digit1<=FOUR; digit2<=ONE; digit3<=ONE; end
      16'd1147: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ONE; digit3<=ONE; end
      16'd1148: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ONE; digit3<=ONE; end
      16'd1149: begin digit0<=NINE; digit1<=FOUR; digit2<=ONE; digit3<=ONE; end
      16'd1150: begin digit0<=ZERO; digit1<=FIVE; digit2<=ONE; digit3<=ONE; end
      16'd1151: begin digit0<=ONE; digit1<=FIVE; digit2<=ONE; digit3<=ONE; end
      16'd1152: begin digit0<=TWO; digit1<=FIVE; digit2<=ONE; digit3<=ONE; end
      16'd1153: begin digit0<=THREE; digit1<=FIVE; digit2<=ONE; digit3<=ONE; end
      16'd1154: begin digit0<=FOUR; digit1<=FIVE; digit2<=ONE; digit3<=ONE; end
      16'd1155: begin digit0<=FIVE; digit1<=FIVE; digit2<=ONE; digit3<=ONE; end
      16'd1156: begin digit0<=SIX; digit1<=FIVE; digit2<=ONE; digit3<=ONE; end
      16'd1157: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ONE; digit3<=ONE; end
      16'd1158: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ONE; digit3<=ONE; end
      16'd1159: begin digit0<=NINE; digit1<=FIVE; digit2<=ONE; digit3<=ONE; end
      16'd1160: begin digit0<=ZERO; digit1<=SIX; digit2<=ONE; digit3<=ONE; end
      16'd1161: begin digit0<=ONE; digit1<=SIX; digit2<=ONE; digit3<=ONE; end
      16'd1162: begin digit0<=TWO; digit1<=SIX; digit2<=ONE; digit3<=ONE; end
      16'd1163: begin digit0<=THREE; digit1<=SIX; digit2<=ONE; digit3<=ONE; end
      16'd1164: begin digit0<=FOUR; digit1<=SIX; digit2<=ONE; digit3<=ONE; end
      16'd1165: begin digit0<=FIVE; digit1<=SIX; digit2<=ONE; digit3<=ONE; end
      16'd1166: begin digit0<=SIX; digit1<=SIX; digit2<=ONE; digit3<=ONE; end
      16'd1167: begin digit0<=SEVEN; digit1<=SIX; digit2<=ONE; digit3<=ONE; end
      16'd1168: begin digit0<=EIGHT; digit1<=SIX; digit2<=ONE; digit3<=ONE; end
      16'd1169: begin digit0<=NINE; digit1<=SIX; digit2<=ONE; digit3<=ONE; end
      16'd1170: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ONE; digit3<=ONE; end
      16'd1171: begin digit0<=ONE; digit1<=SEVEN; digit2<=ONE; digit3<=ONE; end
      16'd1172: begin digit0<=TWO; digit1<=SEVEN; digit2<=ONE; digit3<=ONE; end
      16'd1173: begin digit0<=THREE; digit1<=SEVEN; digit2<=ONE; digit3<=ONE; end
      16'd1174: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ONE; digit3<=ONE; end
      16'd1175: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ONE; digit3<=ONE; end
      16'd1176: begin digit0<=SIX; digit1<=SEVEN; digit2<=ONE; digit3<=ONE; end
      16'd1177: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ONE; digit3<=ONE; end
      16'd1178: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ONE; digit3<=ONE; end
      16'd1179: begin digit0<=NINE; digit1<=SEVEN; digit2<=ONE; digit3<=ONE; end
      16'd1180: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=ONE; end
      16'd1181: begin digit0<=ONE; digit1<=EIGHT; digit2<=ONE; digit3<=ONE; end
      16'd1182: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=ONE; end
      16'd1183: begin digit0<=THREE; digit1<=EIGHT; digit2<=ONE; digit3<=ONE; end
      16'd1184: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ONE; digit3<=ONE; end
      16'd1185: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ONE; digit3<=ONE; end
      16'd1186: begin digit0<=SIX; digit1<=EIGHT; digit2<=ONE; digit3<=ONE; end
      16'd1187: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ONE; digit3<=ONE; end
      16'd1188: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ONE; digit3<=ONE; end
      16'd1189: begin digit0<=NINE; digit1<=EIGHT; digit2<=ONE; digit3<=ONE; end
      16'd1190: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=ONE; end
      16'd1191: begin digit0<=ONE; digit1<=NINE; digit2<=ONE; digit3<=ONE; end
      16'd1192: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=ONE; end
      16'd1193: begin digit0<=THREE; digit1<=NINE; digit2<=ONE; digit3<=ONE; end
      16'd1194: begin digit0<=FOUR; digit1<=NINE; digit2<=ONE; digit3<=ONE; end
      16'd1195: begin digit0<=FIVE; digit1<=NINE; digit2<=ONE; digit3<=ONE; end
      16'd1196: begin digit0<=SIX; digit1<=NINE; digit2<=ONE; digit3<=ONE; end
      16'd1197: begin digit0<=SEVEN; digit1<=NINE; digit2<=ONE; digit3<=ONE; end
      16'd1198: begin digit0<=EIGHT; digit1<=NINE; digit2<=ONE; digit3<=ONE; end
      16'd1199: begin digit0<=NINE; digit1<=NINE; digit2<=ONE; digit3<=ONE; end
	  16'd1200: begin digit0<=ZERO; digit1<=ZERO; digit2<=TWO; digit3<=ONE; end
      16'd1201: begin digit0<=ONE; digit1<=ZERO; digit2<=TWO; digit3<=ONE; end
      16'd1202: begin digit0<=TWO; digit1<=ZERO; digit2<=TWO; digit3<=ONE; end
      16'd1203: begin digit0<=THREE; digit1<=ZERO; digit2<=TWO; digit3<=ONE; end
      16'd1204: begin digit0<=FOUR; digit1<=ZERO; digit2<=TWO; digit3<=ONE; end
      16'd1205: begin digit0<=FIVE; digit1<=ZERO; digit2<=TWO; digit3<=ONE; end
      16'd1206: begin digit0<=SIX; digit1<=ZERO; digit2<=TWO; digit3<=ONE; end
      16'd1207: begin digit0<=SEVEN; digit1<=ZERO; digit2<=TWO; digit3<=ONE; end
      16'd1208: begin digit0<=EIGHT; digit1<=ZERO; digit2<=TWO; digit3<=ONE; end
      16'd1209: begin digit0<=NINE; digit1<=ZERO; digit2<=TWO; digit3<=ONE; end
      16'd1210: begin digit0<=ZERO; digit1<=ONE; digit2<=TWO; digit3<=ONE; end
      16'd1211: begin digit0<=ONE; digit1<=ONE; digit2<=TWO; digit3<=ONE; end
      16'd1212: begin digit0<=TWO; digit1<=ONE; digit2<=TWO; digit3<=ONE; end
      16'd1213: begin digit0<=THREE; digit1<=ONE; digit2<=TWO; digit3<=ONE; end
      16'd1214: begin digit0<=FOUR; digit1<=ONE; digit2<=TWO; digit3<=ONE; end
      16'd1215: begin digit0<=FIVE; digit1<=ONE; digit2<=TWO; digit3<=ONE; end
      16'd1216: begin digit0<=SIX; digit1<=ONE; digit2<=TWO; digit3<=ONE; end
      16'd1217: begin digit0<=SEVEN; digit1<=ONE; digit2<=TWO; digit3<=ONE; end
      16'd1218: begin digit0<=EIGHT; digit1<=ONE; digit2<=TWO; digit3<=ONE; end
      16'd1219: begin digit0<=NINE; digit1<=ONE; digit2<=TWO; digit3<=ONE; end
      16'd1220: begin digit0<=ZERO; digit1<=TWO; digit2<=TWO; digit3<=ONE; end
      16'd1221: begin digit0<=ONE; digit1<=TWO; digit2<=TWO; digit3<=ONE; end
      16'd1222: begin digit0<=TWO; digit1<=TWO; digit2<=TWO; digit3<=ONE; end
      16'd1223: begin digit0<=THREE; digit1<=TWO; digit2<=TWO; digit3<=ONE; end
      16'd1224: begin digit0<=FOUR; digit1<=TWO; digit2<=TWO; digit3<=ONE; end
      16'd1225: begin digit0<=FIVE; digit1<=TWO; digit2<=TWO; digit3<=ONE; end
      16'd1226: begin digit0<=SIX; digit1<=TWO; digit2<=TWO; digit3<=ONE; end
      16'd1227: begin digit0<=SEVEN; digit1<=TWO; digit2<=TWO; digit3<=ONE; end
      16'd1228: begin digit0<=EIGHT; digit1<=TWO; digit2<=TWO; digit3<=ONE; end
      16'd1229: begin digit0<=NINE; digit1<=TWO; digit2<=TWO; digit3<=ONE; end
      16'd1230: begin digit0<=ZERO; digit1<=THREE; digit2<=TWO; digit3<=ONE; end
      16'd1231: begin digit0<=ONE; digit1<=THREE; digit2<=TWO; digit3<=ONE; end
      16'd1232: begin digit0<=TWO; digit1<=THREE; digit2<=TWO; digit3<=ONE; end
      16'd1233: begin digit0<=THREE; digit1<=THREE; digit2<=TWO; digit3<=ONE; end
      16'd1234: begin digit0<=FOUR; digit1<=THREE; digit2<=TWO; digit3<=ONE; end
      16'd1235: begin digit0<=FIVE; digit1<=THREE; digit2<=TWO; digit3<=ONE; end
      16'd1236: begin digit0<=SIX; digit1<=THREE; digit2<=TWO; digit3<=ONE; end
      16'd1237: begin digit0<=SEVEN; digit1<=THREE; digit2<=TWO; digit3<=ONE; end
      16'd1238: begin digit0<=EIGHT; digit1<=THREE; digit2<=TWO; digit3<=ONE; end
      16'd1239: begin digit0<=NINE; digit1<=THREE; digit2<=TWO; digit3<=ONE; end
      16'd1240: begin digit0<=ZERO; digit1<=FOUR; digit2<=TWO; digit3<=ONE; end
      16'd1241: begin digit0<=ONE; digit1<=FOUR; digit2<=TWO; digit3<=ONE; end
      16'd1242: begin digit0<=TWO; digit1<=FOUR; digit2<=TWO; digit3<=ONE; end
      16'd1243: begin digit0<=THREE; digit1<=FOUR; digit2<=TWO; digit3<=ONE; end
      16'd1244: begin digit0<=FOUR; digit1<=FOUR; digit2<=TWO; digit3<=ONE; end
      16'd1245: begin digit0<=FIVE; digit1<=FOUR; digit2<=TWO; digit3<=ONE; end
      16'd1246: begin digit0<=SIX; digit1<=FOUR; digit2<=TWO; digit3<=ONE; end
      16'd1247: begin digit0<=SEVEN; digit1<=FOUR; digit2<=TWO; digit3<=ONE; end
      16'd1248: begin digit0<=EIGHT; digit1<=FOUR; digit2<=TWO; digit3<=ONE; end
      16'd1249: begin digit0<=NINE; digit1<=FOUR; digit2<=TWO; digit3<=ONE; end
      16'd1250: begin digit0<=ZERO; digit1<=FIVE; digit2<=TWO; digit3<=ONE; end
      16'd1251: begin digit0<=ONE; digit1<=FIVE; digit2<=TWO; digit3<=ONE; end
      16'd1252: begin digit0<=TWO; digit1<=FIVE; digit2<=TWO; digit3<=ONE; end
      16'd1253: begin digit0<=THREE; digit1<=FIVE; digit2<=TWO; digit3<=ONE; end
      16'd1254: begin digit0<=FOUR; digit1<=FIVE; digit2<=TWO; digit3<=ONE; end
      16'd1255: begin digit0<=FIVE; digit1<=FIVE; digit2<=TWO; digit3<=ONE; end
      16'd1256: begin digit0<=SIX; digit1<=FIVE; digit2<=TWO; digit3<=ONE; end
      16'd1257: begin digit0<=SEVEN; digit1<=FIVE; digit2<=TWO; digit3<=ONE; end
      16'd1258: begin digit0<=EIGHT; digit1<=FIVE; digit2<=TWO; digit3<=ONE; end
      16'd1259: begin digit0<=NINE; digit1<=FIVE; digit2<=TWO; digit3<=ONE; end
      16'd1260: begin digit0<=ZERO; digit1<=SIX; digit2<=TWO; digit3<=ONE; end
      16'd1261: begin digit0<=ONE; digit1<=SIX; digit2<=TWO; digit3<=ONE; end
      16'd1262: begin digit0<=TWO; digit1<=SIX; digit2<=TWO; digit3<=ONE; end
      16'd1263: begin digit0<=THREE; digit1<=SIX; digit2<=TWO; digit3<=ONE; end
      16'd1264: begin digit0<=FOUR; digit1<=SIX; digit2<=TWO; digit3<=ONE; end
      16'd1265: begin digit0<=FIVE; digit1<=SIX; digit2<=TWO; digit3<=ONE; end
      16'd1266: begin digit0<=SIX; digit1<=SIX; digit2<=TWO; digit3<=ONE; end
      16'd1267: begin digit0<=SEVEN; digit1<=SIX; digit2<=TWO; digit3<=ONE; end
      16'd1268: begin digit0<=EIGHT; digit1<=SIX; digit2<=TWO; digit3<=ONE; end
      16'd1269: begin digit0<=NINE; digit1<=SIX; digit2<=TWO; digit3<=ONE; end
      16'd1270: begin digit0<=ZERO; digit1<=SEVEN; digit2<=TWO; digit3<=ONE; end
      16'd1271: begin digit0<=ONE; digit1<=SEVEN; digit2<=TWO; digit3<=ONE; end
      16'd1272: begin digit0<=TWO; digit1<=SEVEN; digit2<=TWO; digit3<=ONE; end
      16'd1273: begin digit0<=THREE; digit1<=SEVEN; digit2<=TWO; digit3<=ONE; end
      16'd1274: begin digit0<=FOUR; digit1<=SEVEN; digit2<=TWO; digit3<=ONE; end
      16'd1275: begin digit0<=FIVE; digit1<=SEVEN; digit2<=TWO; digit3<=ONE; end
      16'd1276: begin digit0<=SIX; digit1<=SEVEN; digit2<=TWO; digit3<=ONE; end
      16'd1277: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=TWO; digit3<=ONE; end
      16'd1278: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=TWO; digit3<=ONE; end
      16'd1279: begin digit0<=NINE; digit1<=SEVEN; digit2<=TWO; digit3<=ONE; end
      16'd1280: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=ONE; end
      16'd1281: begin digit0<=ONE; digit1<=EIGHT; digit2<=TWO; digit3<=ONE; end
      16'd1282: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=ONE; end
      16'd1283: begin digit0<=THREE; digit1<=EIGHT; digit2<=TWO; digit3<=ONE; end
      16'd1284: begin digit0<=FOUR; digit1<=EIGHT; digit2<=TWO; digit3<=ONE; end
      16'd1285: begin digit0<=FIVE; digit1<=EIGHT; digit2<=TWO; digit3<=ONE; end
      16'd1286: begin digit0<=SIX; digit1<=EIGHT; digit2<=TWO; digit3<=ONE; end
      16'd1287: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=TWO; digit3<=ONE; end
      16'd1288: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=TWO; digit3<=ONE; end
      16'd1289: begin digit0<=NINE; digit1<=EIGHT; digit2<=TWO; digit3<=ONE; end
      16'd1290: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=ONE; end
      16'd1291: begin digit0<=ONE; digit1<=NINE; digit2<=TWO; digit3<=ONE; end
      16'd1292: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=ONE; end
      16'd1293: begin digit0<=THREE; digit1<=NINE; digit2<=TWO; digit3<=ONE; end
      16'd1294: begin digit0<=FOUR; digit1<=NINE; digit2<=TWO; digit3<=ONE; end
      16'd1295: begin digit0<=FIVE; digit1<=NINE; digit2<=TWO; digit3<=ONE; end
      16'd1296: begin digit0<=SIX; digit1<=NINE; digit2<=TWO; digit3<=ONE; end
      16'd1297: begin digit0<=SEVEN; digit1<=NINE; digit2<=TWO; digit3<=ONE; end
      16'd1298: begin digit0<=EIGHT; digit1<=NINE; digit2<=TWO; digit3<=ONE; end
      16'd1299: begin digit0<=NINE; digit1<=NINE; digit2<=TWO; digit3<=ONE; end
	  16'd1300: begin digit0<=ZERO; digit1<=ZERO; digit2<=THREE; digit3<=ONE; end
      16'd1301: begin digit0<=ONE; digit1<=ZERO; digit2<=THREE; digit3<=ONE; end
      16'd1302: begin digit0<=TWO; digit1<=ZERO; digit2<=THREE; digit3<=ONE; end
      16'd1303: begin digit0<=THREE; digit1<=ZERO; digit2<=THREE; digit3<=ONE; end
      16'd1304: begin digit0<=FOUR; digit1<=ZERO; digit2<=THREE; digit3<=ONE; end
      16'd1305: begin digit0<=FIVE; digit1<=ZERO; digit2<=THREE; digit3<=ONE; end
      16'd1306: begin digit0<=SIX; digit1<=ZERO; digit2<=THREE; digit3<=ONE; end
      16'd1307: begin digit0<=SEVEN; digit1<=ZERO; digit2<=THREE; digit3<=ONE; end
      16'd1308: begin digit0<=EIGHT; digit1<=ZERO; digit2<=THREE; digit3<=ONE; end
      16'd1309: begin digit0<=NINE; digit1<=ZERO; digit2<=THREE; digit3<=ONE; end
      16'd1310: begin digit0<=ZERO; digit1<=ONE; digit2<=THREE; digit3<=ONE; end
      16'd1311: begin digit0<=ONE; digit1<=ONE; digit2<=THREE; digit3<=ONE; end
      16'd1312: begin digit0<=TWO; digit1<=ONE; digit2<=THREE; digit3<=ONE; end
      16'd1313: begin digit0<=THREE; digit1<=ONE; digit2<=THREE; digit3<=ONE; end
      16'd1314: begin digit0<=FOUR; digit1<=ONE; digit2<=THREE; digit3<=ONE; end
      16'd1315: begin digit0<=FIVE; digit1<=ONE; digit2<=THREE; digit3<=ONE; end
      16'd1316: begin digit0<=SIX; digit1<=ONE; digit2<=THREE; digit3<=ONE; end
      16'd1317: begin digit0<=SEVEN; digit1<=ONE; digit2<=THREE; digit3<=ONE; end
      16'd1318: begin digit0<=EIGHT; digit1<=ONE; digit2<=THREE; digit3<=ONE; end
      16'd1319: begin digit0<=NINE; digit1<=ONE; digit2<=THREE; digit3<=ONE; end
      16'd1320: begin digit0<=ZERO; digit1<=TWO; digit2<=THREE; digit3<=ONE; end
      16'd1321: begin digit0<=ONE; digit1<=TWO; digit2<=THREE; digit3<=ONE; end
      16'd1322: begin digit0<=TWO; digit1<=TWO; digit2<=THREE; digit3<=ONE; end
      16'd1323: begin digit0<=THREE; digit1<=TWO; digit2<=THREE; digit3<=ONE; end
      16'd1324: begin digit0<=FOUR; digit1<=TWO; digit2<=THREE; digit3<=ONE; end
      16'd1325: begin digit0<=FIVE; digit1<=TWO; digit2<=THREE; digit3<=ONE; end
      16'd1326: begin digit0<=SIX; digit1<=TWO; digit2<=THREE; digit3<=ONE; end
      16'd1327: begin digit0<=SEVEN; digit1<=TWO; digit2<=THREE; digit3<=ONE; end
      16'd1328: begin digit0<=EIGHT; digit1<=TWO; digit2<=THREE; digit3<=ONE; end
      16'd1329: begin digit0<=NINE; digit1<=TWO; digit2<=THREE; digit3<=ONE; end
      16'd1330: begin digit0<=ZERO; digit1<=THREE; digit2<=THREE; digit3<=ONE; end
      16'd1331: begin digit0<=ONE; digit1<=THREE; digit2<=THREE; digit3<=ONE; end
      16'd1332: begin digit0<=TWO; digit1<=THREE; digit2<=THREE; digit3<=ONE; end
      16'd1333: begin digit0<=THREE; digit1<=THREE; digit2<=THREE; digit3<=ONE; end
      16'd1334: begin digit0<=FOUR; digit1<=THREE; digit2<=THREE; digit3<=ONE; end
      16'd1335: begin digit0<=FIVE; digit1<=THREE; digit2<=THREE; digit3<=ONE; end
      16'd1336: begin digit0<=SIX; digit1<=THREE; digit2<=THREE; digit3<=ONE; end
      16'd1337: begin digit0<=SEVEN; digit1<=THREE; digit2<=THREE; digit3<=ONE; end
      16'd1338: begin digit0<=EIGHT; digit1<=THREE; digit2<=THREE; digit3<=ONE; end
      16'd1339: begin digit0<=NINE; digit1<=THREE; digit2<=THREE; digit3<=ONE; end
      16'd1340: begin digit0<=ZERO; digit1<=FOUR; digit2<=THREE; digit3<=ONE; end
      16'd1341: begin digit0<=ONE; digit1<=FOUR; digit2<=THREE; digit3<=ONE; end
      16'd1342: begin digit0<=TWO; digit1<=FOUR; digit2<=THREE; digit3<=ONE; end
      16'd1343: begin digit0<=THREE; digit1<=FOUR; digit2<=THREE; digit3<=ONE; end
      16'd1344: begin digit0<=FOUR; digit1<=FOUR; digit2<=THREE; digit3<=ONE; end
      16'd1345: begin digit0<=FIVE; digit1<=FOUR; digit2<=THREE; digit3<=ONE; end
      16'd1346: begin digit0<=SIX; digit1<=FOUR; digit2<=THREE; digit3<=ONE; end
      16'd1347: begin digit0<=SEVEN; digit1<=FOUR; digit2<=THREE; digit3<=ONE; end
      16'd1348: begin digit0<=EIGHT; digit1<=FOUR; digit2<=THREE; digit3<=ONE; end
      16'd1349: begin digit0<=NINE; digit1<=FOUR; digit2<=THREE; digit3<=ONE; end
      16'd1350: begin digit0<=ZERO; digit1<=FIVE; digit2<=THREE; digit3<=ONE; end
      16'd1351: begin digit0<=ONE; digit1<=FIVE; digit2<=THREE; digit3<=ONE; end
      16'd1352: begin digit0<=TWO; digit1<=FIVE; digit2<=THREE; digit3<=ONE; end
      16'd1353: begin digit0<=THREE; digit1<=FIVE; digit2<=THREE; digit3<=ONE; end
      16'd1354: begin digit0<=FOUR; digit1<=FIVE; digit2<=THREE; digit3<=ONE; end
      16'd1355: begin digit0<=FIVE; digit1<=FIVE; digit2<=THREE; digit3<=ONE; end
      16'd1356: begin digit0<=SIX; digit1<=FIVE; digit2<=THREE; digit3<=ONE; end
      16'd1357: begin digit0<=SEVEN; digit1<=FIVE; digit2<=THREE; digit3<=ONE; end
      16'd1358: begin digit0<=EIGHT; digit1<=FIVE; digit2<=THREE; digit3<=ONE; end
      16'd1359: begin digit0<=NINE; digit1<=FIVE; digit2<=THREE; digit3<=ONE; end
      16'd1360: begin digit0<=ZERO; digit1<=SIX; digit2<=THREE; digit3<=ONE; end
      16'd1361: begin digit0<=ONE; digit1<=SIX; digit2<=THREE; digit3<=ONE; end
      16'd1362: begin digit0<=TWO; digit1<=SIX; digit2<=THREE; digit3<=ONE; end
      16'd1363: begin digit0<=THREE; digit1<=SIX; digit2<=THREE; digit3<=ONE; end
      16'd1364: begin digit0<=FOUR; digit1<=SIX; digit2<=THREE; digit3<=ONE; end
      16'd1365: begin digit0<=FIVE; digit1<=SIX; digit2<=THREE; digit3<=ONE; end
      16'd1366: begin digit0<=SIX; digit1<=SIX; digit2<=THREE; digit3<=ONE; end
      16'd1367: begin digit0<=SEVEN; digit1<=SIX; digit2<=THREE; digit3<=ONE; end
      16'd1368: begin digit0<=EIGHT; digit1<=SIX; digit2<=THREE; digit3<=ONE; end
      16'd1369: begin digit0<=NINE; digit1<=SIX; digit2<=THREE; digit3<=ONE; end
      16'd1370: begin digit0<=ZERO; digit1<=SEVEN; digit2<=THREE; digit3<=ONE; end
      16'd1371: begin digit0<=ONE; digit1<=SEVEN; digit2<=THREE; digit3<=ONE; end
      16'd1372: begin digit0<=TWO; digit1<=SEVEN; digit2<=THREE; digit3<=ONE; end
      16'd1373: begin digit0<=THREE; digit1<=SEVEN; digit2<=THREE; digit3<=ONE; end
      16'd1374: begin digit0<=FOUR; digit1<=SEVEN; digit2<=THREE; digit3<=ONE; end
      16'd1375: begin digit0<=FIVE; digit1<=SEVEN; digit2<=THREE; digit3<=ONE; end
      16'd1376: begin digit0<=SIX; digit1<=SEVEN; digit2<=THREE; digit3<=ONE; end
      16'd1377: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=THREE; digit3<=ONE; end
      16'd1378: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=THREE; digit3<=ONE; end
      16'd1379: begin digit0<=NINE; digit1<=SEVEN; digit2<=THREE; digit3<=ONE; end
      16'd1380: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=ONE; end
      16'd1381: begin digit0<=ONE; digit1<=EIGHT; digit2<=THREE; digit3<=ONE; end
      16'd1382: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=ONE; end
      16'd1383: begin digit0<=THREE; digit1<=EIGHT; digit2<=THREE; digit3<=ONE; end
      16'd1384: begin digit0<=FOUR; digit1<=EIGHT; digit2<=THREE; digit3<=ONE; end
      16'd1385: begin digit0<=FIVE; digit1<=EIGHT; digit2<=THREE; digit3<=ONE; end
      16'd1386: begin digit0<=SIX; digit1<=EIGHT; digit2<=THREE; digit3<=ONE; end
      16'd1387: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=THREE; digit3<=ONE; end
      16'd1388: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=THREE; digit3<=ONE; end
      16'd1389: begin digit0<=NINE; digit1<=EIGHT; digit2<=THREE; digit3<=ONE; end
      16'd1390: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=ONE; end
      16'd1391: begin digit0<=ONE; digit1<=NINE; digit2<=THREE; digit3<=ONE; end
      16'd1392: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=ONE; end
      16'd1393: begin digit0<=THREE; digit1<=NINE; digit2<=THREE; digit3<=ONE; end
      16'd1394: begin digit0<=FOUR; digit1<=NINE; digit2<=THREE; digit3<=ONE; end
      16'd1395: begin digit0<=FIVE; digit1<=NINE; digit2<=THREE; digit3<=ONE; end
      16'd1396: begin digit0<=SIX; digit1<=NINE; digit2<=THREE; digit3<=ONE; end
      16'd1397: begin digit0<=SEVEN; digit1<=NINE; digit2<=THREE; digit3<=ONE; end
      16'd1398: begin digit0<=EIGHT; digit1<=NINE; digit2<=THREE; digit3<=ONE; end
      16'd1399: begin digit0<=NINE; digit1<=NINE; digit2<=THREE; digit3<=ONE; end
	  16'd1400: begin digit0<=ZERO; digit1<=ZERO; digit2<=FOUR; digit3<=ONE; end
      16'd1401: begin digit0<=ONE; digit1<=ZERO; digit2<=FOUR; digit3<=ONE; end
      16'd1402: begin digit0<=TWO; digit1<=ZERO; digit2<=FOUR; digit3<=ONE; end
      16'd1403: begin digit0<=THREE; digit1<=ZERO; digit2<=FOUR; digit3<=ONE; end
      16'd1404: begin digit0<=FOUR; digit1<=ZERO; digit2<=FOUR; digit3<=ONE; end
      16'd1405: begin digit0<=FIVE; digit1<=ZERO; digit2<=FOUR; digit3<=ONE; end
      16'd1406: begin digit0<=SIX; digit1<=ZERO; digit2<=FOUR; digit3<=ONE; end
      16'd1407: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FOUR; digit3<=ONE; end
      16'd1408: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FOUR; digit3<=ONE; end
      16'd1409: begin digit0<=NINE; digit1<=ZERO; digit2<=FOUR; digit3<=ONE; end
      16'd1410: begin digit0<=ZERO; digit1<=ONE; digit2<=FOUR; digit3<=ONE; end
      16'd1411: begin digit0<=ONE; digit1<=ONE; digit2<=FOUR; digit3<=ONE; end
      16'd1412: begin digit0<=TWO; digit1<=ONE; digit2<=FOUR; digit3<=ONE; end
      16'd1413: begin digit0<=THREE; digit1<=ONE; digit2<=FOUR; digit3<=ONE; end
      16'd1414: begin digit0<=FOUR; digit1<=ONE; digit2<=FOUR; digit3<=ONE; end
      16'd1415: begin digit0<=FIVE; digit1<=ONE; digit2<=FOUR; digit3<=ONE; end
      16'd1416: begin digit0<=SIX; digit1<=ONE; digit2<=FOUR; digit3<=ONE; end
      16'd1417: begin digit0<=SEVEN; digit1<=ONE; digit2<=FOUR; digit3<=ONE; end
      16'd1418: begin digit0<=EIGHT; digit1<=ONE; digit2<=FOUR; digit3<=ONE; end
      16'd1419: begin digit0<=NINE; digit1<=ONE; digit2<=FOUR; digit3<=ONE; end
      16'd1420: begin digit0<=ZERO; digit1<=TWO; digit2<=FOUR; digit3<=ONE; end
      16'd1421: begin digit0<=ONE; digit1<=TWO; digit2<=FOUR; digit3<=ONE; end
      16'd1422: begin digit0<=TWO; digit1<=TWO; digit2<=FOUR; digit3<=ONE; end
      16'd1423: begin digit0<=THREE; digit1<=TWO; digit2<=FOUR; digit3<=ONE; end
      16'd1424: begin digit0<=FOUR; digit1<=TWO; digit2<=FOUR; digit3<=ONE; end
      16'd1425: begin digit0<=FIVE; digit1<=TWO; digit2<=FOUR; digit3<=ONE; end
      16'd1426: begin digit0<=SIX; digit1<=TWO; digit2<=FOUR; digit3<=ONE; end
      16'd1427: begin digit0<=SEVEN; digit1<=TWO; digit2<=FOUR; digit3<=ONE; end
      16'd1428: begin digit0<=EIGHT; digit1<=TWO; digit2<=FOUR; digit3<=ONE; end
      16'd1429: begin digit0<=NINE; digit1<=TWO; digit2<=FOUR; digit3<=ONE; end
      16'd1430: begin digit0<=ZERO; digit1<=THREE; digit2<=FOUR; digit3<=ONE; end
      16'd1431: begin digit0<=ONE; digit1<=THREE; digit2<=FOUR; digit3<=ONE; end
      16'd1432: begin digit0<=TWO; digit1<=THREE; digit2<=FOUR; digit3<=ONE; end
      16'd1433: begin digit0<=THREE; digit1<=THREE; digit2<=FOUR; digit3<=ONE; end
      16'd1434: begin digit0<=FOUR; digit1<=THREE; digit2<=FOUR; digit3<=ONE; end
      16'd1435: begin digit0<=FIVE; digit1<=THREE; digit2<=FOUR; digit3<=ONE; end
      16'd1436: begin digit0<=SIX; digit1<=THREE; digit2<=FOUR; digit3<=ONE; end
      16'd1437: begin digit0<=SEVEN; digit1<=THREE; digit2<=FOUR; digit3<=ONE; end
      16'd1438: begin digit0<=EIGHT; digit1<=THREE; digit2<=FOUR; digit3<=ONE; end
      16'd1439: begin digit0<=NINE; digit1<=THREE; digit2<=FOUR; digit3<=ONE; end
      16'd1440: begin digit0<=ZERO; digit1<=FOUR; digit2<=FOUR; digit3<=ONE; end
      16'd1441: begin digit0<=ONE; digit1<=FOUR; digit2<=FOUR; digit3<=ONE; end
      16'd1442: begin digit0<=TWO; digit1<=FOUR; digit2<=FOUR; digit3<=ONE; end
      16'd1443: begin digit0<=THREE; digit1<=FOUR; digit2<=FOUR; digit3<=ONE; end
      16'd1444: begin digit0<=FOUR; digit1<=FOUR; digit2<=FOUR; digit3<=ONE; end
      16'd1445: begin digit0<=FIVE; digit1<=FOUR; digit2<=FOUR; digit3<=ONE; end
      16'd1446: begin digit0<=SIX; digit1<=FOUR; digit2<=FOUR; digit3<=ONE; end
      16'd1447: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FOUR; digit3<=ONE; end
      16'd1448: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FOUR; digit3<=ONE; end
      16'd1449: begin digit0<=NINE; digit1<=FOUR; digit2<=FOUR; digit3<=ONE; end
      16'd1450: begin digit0<=ZERO; digit1<=FIVE; digit2<=FOUR; digit3<=ONE; end
      16'd1451: begin digit0<=ONE; digit1<=FIVE; digit2<=FOUR; digit3<=ONE; end
      16'd1452: begin digit0<=TWO; digit1<=FIVE; digit2<=FOUR; digit3<=ONE; end
      16'd1453: begin digit0<=THREE; digit1<=FIVE; digit2<=FOUR; digit3<=ONE; end
      16'd1454: begin digit0<=FOUR; digit1<=FIVE; digit2<=FOUR; digit3<=ONE; end
      16'd1455: begin digit0<=FIVE; digit1<=FIVE; digit2<=FOUR; digit3<=ONE; end
      16'd1456: begin digit0<=SIX; digit1<=FIVE; digit2<=FOUR; digit3<=ONE; end
      16'd1457: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FOUR; digit3<=ONE; end
      16'd1458: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FOUR; digit3<=ONE; end
      16'd1459: begin digit0<=NINE; digit1<=FIVE; digit2<=FOUR; digit3<=ONE; end
      16'd1460: begin digit0<=ZERO; digit1<=SIX; digit2<=FOUR; digit3<=ONE; end
      16'd1461: begin digit0<=ONE; digit1<=SIX; digit2<=FOUR; digit3<=ONE; end
      16'd1462: begin digit0<=TWO; digit1<=SIX; digit2<=FOUR; digit3<=ONE; end
      16'd1463: begin digit0<=THREE; digit1<=SIX; digit2<=FOUR; digit3<=ONE; end
      16'd1464: begin digit0<=FOUR; digit1<=SIX; digit2<=FOUR; digit3<=ONE; end
      16'd1465: begin digit0<=FIVE; digit1<=SIX; digit2<=FOUR; digit3<=ONE; end
      16'd1466: begin digit0<=SIX; digit1<=SIX; digit2<=FOUR; digit3<=ONE; end
      16'd1467: begin digit0<=SEVEN; digit1<=SIX; digit2<=FOUR; digit3<=ONE; end
      16'd1468: begin digit0<=EIGHT; digit1<=SIX; digit2<=FOUR; digit3<=ONE; end
      16'd1469: begin digit0<=NINE; digit1<=SIX; digit2<=FOUR; digit3<=ONE; end
      16'd1470: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FOUR; digit3<=ONE; end
      16'd1471: begin digit0<=ONE; digit1<=SEVEN; digit2<=FOUR; digit3<=ONE; end
      16'd1472: begin digit0<=TWO; digit1<=SEVEN; digit2<=FOUR; digit3<=ONE; end
      16'd1473: begin digit0<=THREE; digit1<=SEVEN; digit2<=FOUR; digit3<=ONE; end
      16'd1474: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FOUR; digit3<=ONE; end
      16'd1475: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FOUR; digit3<=ONE; end
      16'd1476: begin digit0<=SIX; digit1<=SEVEN; digit2<=FOUR; digit3<=ONE; end
      16'd1477: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FOUR; digit3<=ONE; end
      16'd1478: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FOUR; digit3<=ONE; end
      16'd1479: begin digit0<=NINE; digit1<=SEVEN; digit2<=FOUR; digit3<=ONE; end
      16'd1480: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=ONE; end
      16'd1481: begin digit0<=ONE; digit1<=EIGHT; digit2<=FOUR; digit3<=ONE; end
      16'd1482: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=ONE; end
      16'd1483: begin digit0<=THREE; digit1<=EIGHT; digit2<=FOUR; digit3<=ONE; end
      16'd1484: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FOUR; digit3<=ONE; end
      16'd1485: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FOUR; digit3<=ONE; end
      16'd1486: begin digit0<=SIX; digit1<=EIGHT; digit2<=FOUR; digit3<=ONE; end
      16'd1487: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FOUR; digit3<=ONE; end
      16'd1488: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FOUR; digit3<=ONE; end
      16'd1489: begin digit0<=NINE; digit1<=EIGHT; digit2<=FOUR; digit3<=ONE; end
      16'd1490: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=ONE; end
      16'd1491: begin digit0<=ONE; digit1<=NINE; digit2<=FOUR; digit3<=ONE; end
      16'd1492: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=ONE; end
      16'd1493: begin digit0<=THREE; digit1<=NINE; digit2<=FOUR; digit3<=ONE; end
      16'd1494: begin digit0<=FOUR; digit1<=NINE; digit2<=FOUR; digit3<=ONE; end
      16'd1495: begin digit0<=FIVE; digit1<=NINE; digit2<=FOUR; digit3<=ONE; end
      16'd1496: begin digit0<=SIX; digit1<=NINE; digit2<=FOUR; digit3<=ONE; end
      16'd1497: begin digit0<=SEVEN; digit1<=NINE; digit2<=FOUR; digit3<=ONE; end
      16'd1498: begin digit0<=EIGHT; digit1<=NINE; digit2<=FOUR; digit3<=ONE; end
      16'd1499: begin digit0<=NINE; digit1<=NINE; digit2<=FOUR; digit3<=ONE; end
	  16'd1500: begin digit0<=ZERO; digit1<=ZERO; digit2<=FIVE; digit3<=ONE; end
      16'd1501: begin digit0<=ONE; digit1<=ZERO; digit2<=FIVE; digit3<=ONE; end
      16'd1502: begin digit0<=TWO; digit1<=ZERO; digit2<=FIVE; digit3<=ONE; end
      16'd1503: begin digit0<=THREE; digit1<=ZERO; digit2<=FIVE; digit3<=ONE; end
      16'd1504: begin digit0<=FOUR; digit1<=ZERO; digit2<=FIVE; digit3<=ONE; end
      16'd1505: begin digit0<=FIVE; digit1<=ZERO; digit2<=FIVE; digit3<=ONE; end
      16'd1506: begin digit0<=SIX; digit1<=ZERO; digit2<=FIVE; digit3<=ONE; end
      16'd1507: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FIVE; digit3<=ONE; end
      16'd1508: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FIVE; digit3<=ONE; end
      16'd1509: begin digit0<=NINE; digit1<=ZERO; digit2<=FIVE; digit3<=ONE; end
      16'd1510: begin digit0<=ZERO; digit1<=ONE; digit2<=FIVE; digit3<=ONE; end
      16'd1511: begin digit0<=ONE; digit1<=ONE; digit2<=FIVE; digit3<=ONE; end
      16'd1512: begin digit0<=TWO; digit1<=ONE; digit2<=FIVE; digit3<=ONE; end
      16'd1513: begin digit0<=THREE; digit1<=ONE; digit2<=FIVE; digit3<=ONE; end
      16'd1514: begin digit0<=FOUR; digit1<=ONE; digit2<=FIVE; digit3<=ONE; end
      16'd1515: begin digit0<=FIVE; digit1<=ONE; digit2<=FIVE; digit3<=ONE; end
      16'd1516: begin digit0<=SIX; digit1<=ONE; digit2<=FIVE; digit3<=ONE; end
      16'd1517: begin digit0<=SEVEN; digit1<=ONE; digit2<=FIVE; digit3<=ONE; end
      16'd1518: begin digit0<=EIGHT; digit1<=ONE; digit2<=FIVE; digit3<=ONE; end
      16'd1519: begin digit0<=NINE; digit1<=ONE; digit2<=FIVE; digit3<=ONE; end
      16'd1520: begin digit0<=ZERO; digit1<=TWO; digit2<=FIVE; digit3<=ONE; end
      16'd1521: begin digit0<=ONE; digit1<=TWO; digit2<=FIVE; digit3<=ONE; end
      16'd1522: begin digit0<=TWO; digit1<=TWO; digit2<=FIVE; digit3<=ONE; end
      16'd1523: begin digit0<=THREE; digit1<=TWO; digit2<=FIVE; digit3<=ONE; end
      16'd1524: begin digit0<=FOUR; digit1<=TWO; digit2<=FIVE; digit3<=ONE; end
      16'd1525: begin digit0<=FIVE; digit1<=TWO; digit2<=FIVE; digit3<=ONE; end
      16'd1526: begin digit0<=SIX; digit1<=TWO; digit2<=FIVE; digit3<=ONE; end
      16'd1527: begin digit0<=SEVEN; digit1<=TWO; digit2<=FIVE; digit3<=ONE; end
      16'd1528: begin digit0<=EIGHT; digit1<=TWO; digit2<=FIVE; digit3<=ONE; end
      16'd1529: begin digit0<=NINE; digit1<=TWO; digit2<=FIVE; digit3<=ONE; end
      16'd1530: begin digit0<=ZERO; digit1<=THREE; digit2<=FIVE; digit3<=ONE; end
      16'd1531: begin digit0<=ONE; digit1<=THREE; digit2<=FIVE; digit3<=ONE; end
      16'd1532: begin digit0<=TWO; digit1<=THREE; digit2<=FIVE; digit3<=ONE; end
      16'd1533: begin digit0<=THREE; digit1<=THREE; digit2<=FIVE; digit3<=ONE; end
      16'd1534: begin digit0<=FOUR; digit1<=THREE; digit2<=FIVE; digit3<=ONE; end
      16'd1535: begin digit0<=FIVE; digit1<=THREE; digit2<=FIVE; digit3<=ONE; end
      16'd1536: begin digit0<=SIX; digit1<=THREE; digit2<=FIVE; digit3<=ONE; end
      16'd1537: begin digit0<=SEVEN; digit1<=THREE; digit2<=FIVE; digit3<=ONE; end
      16'd1538: begin digit0<=EIGHT; digit1<=THREE; digit2<=FIVE; digit3<=ONE; end
      16'd1539: begin digit0<=NINE; digit1<=THREE; digit2<=FIVE; digit3<=ONE; end
      16'd1540: begin digit0<=ZERO; digit1<=FOUR; digit2<=FIVE; digit3<=ONE; end
      16'd1541: begin digit0<=ONE; digit1<=FOUR; digit2<=FIVE; digit3<=ONE; end
      16'd1542: begin digit0<=TWO; digit1<=FOUR; digit2<=FIVE; digit3<=ONE; end
      16'd1543: begin digit0<=THREE; digit1<=FOUR; digit2<=FIVE; digit3<=ONE; end
      16'd1544: begin digit0<=FOUR; digit1<=FOUR; digit2<=FIVE; digit3<=ONE; end
      16'd1545: begin digit0<=FIVE; digit1<=FOUR; digit2<=FIVE; digit3<=ONE; end
      16'd1546: begin digit0<=SIX; digit1<=FOUR; digit2<=FIVE; digit3<=ONE; end
      16'd1547: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FIVE; digit3<=ONE; end
      16'd1548: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FIVE; digit3<=ONE; end
      16'd1549: begin digit0<=NINE; digit1<=FOUR; digit2<=FIVE; digit3<=ONE; end
      16'd1550: begin digit0<=ZERO; digit1<=FIVE; digit2<=FIVE; digit3<=ONE; end
      16'd1551: begin digit0<=ONE; digit1<=FIVE; digit2<=FIVE; digit3<=ONE; end
      16'd1552: begin digit0<=TWO; digit1<=FIVE; digit2<=FIVE; digit3<=ONE; end
      16'd1553: begin digit0<=THREE; digit1<=FIVE; digit2<=FIVE; digit3<=ONE; end
      16'd1554: begin digit0<=FOUR; digit1<=FIVE; digit2<=FIVE; digit3<=ONE; end
      16'd1555: begin digit0<=FIVE; digit1<=FIVE; digit2<=FIVE; digit3<=ONE; end
      16'd1556: begin digit0<=SIX; digit1<=FIVE; digit2<=FIVE; digit3<=ONE; end
      16'd1557: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FIVE; digit3<=ONE; end
      16'd1558: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FIVE; digit3<=ONE; end
      16'd1559: begin digit0<=NINE; digit1<=FIVE; digit2<=FIVE; digit3<=ONE; end
      16'd1560: begin digit0<=ZERO; digit1<=SIX; digit2<=FIVE; digit3<=ONE; end
      16'd1561: begin digit0<=ONE; digit1<=SIX; digit2<=FIVE; digit3<=ONE; end
      16'd1562: begin digit0<=TWO; digit1<=SIX; digit2<=FIVE; digit3<=ONE; end
      16'd1563: begin digit0<=THREE; digit1<=SIX; digit2<=FIVE; digit3<=ONE; end
      16'd1564: begin digit0<=FOUR; digit1<=SIX; digit2<=FIVE; digit3<=ONE; end
      16'd1565: begin digit0<=FIVE; digit1<=SIX; digit2<=FIVE; digit3<=ONE; end
      16'd1566: begin digit0<=SIX; digit1<=SIX; digit2<=FIVE; digit3<=ONE; end
      16'd1567: begin digit0<=SEVEN; digit1<=SIX; digit2<=FIVE; digit3<=ONE; end
      16'd1568: begin digit0<=EIGHT; digit1<=SIX; digit2<=FIVE; digit3<=ONE; end
      16'd1569: begin digit0<=NINE; digit1<=SIX; digit2<=FIVE; digit3<=ONE; end
      16'd1570: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FIVE; digit3<=ONE; end
      16'd1571: begin digit0<=ONE; digit1<=SEVEN; digit2<=FIVE; digit3<=ONE; end
      16'd1572: begin digit0<=TWO; digit1<=SEVEN; digit2<=FIVE; digit3<=ONE; end
      16'd1573: begin digit0<=THREE; digit1<=SEVEN; digit2<=FIVE; digit3<=ONE; end
      16'd1574: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FIVE; digit3<=ONE; end
      16'd1575: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FIVE; digit3<=ONE; end
      16'd1576: begin digit0<=SIX; digit1<=SEVEN; digit2<=FIVE; digit3<=ONE; end
      16'd1577: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FIVE; digit3<=ONE; end
      16'd1578: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FIVE; digit3<=ONE; end
      16'd1579: begin digit0<=NINE; digit1<=SEVEN; digit2<=FIVE; digit3<=ONE; end
      16'd1580: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=ONE; end
      16'd1581: begin digit0<=ONE; digit1<=EIGHT; digit2<=FIVE; digit3<=ONE; end
      16'd1582: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=ONE; end
      16'd1583: begin digit0<=THREE; digit1<=EIGHT; digit2<=FIVE; digit3<=ONE; end
      16'd1584: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FIVE; digit3<=ONE; end
      16'd1585: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FIVE; digit3<=ONE; end
      16'd1586: begin digit0<=SIX; digit1<=EIGHT; digit2<=FIVE; digit3<=ONE; end
      16'd1587: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FIVE; digit3<=ONE; end
      16'd1588: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FIVE; digit3<=ONE; end
      16'd1589: begin digit0<=NINE; digit1<=EIGHT; digit2<=FIVE; digit3<=ONE; end
      16'd1590: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=ONE; end
      16'd1591: begin digit0<=ONE; digit1<=NINE; digit2<=FIVE; digit3<=ONE; end
      16'd1592: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=ONE; end
      16'd1593: begin digit0<=THREE; digit1<=NINE; digit2<=FIVE; digit3<=ONE; end
      16'd1594: begin digit0<=FOUR; digit1<=NINE; digit2<=FIVE; digit3<=ONE; end
      16'd1595: begin digit0<=FIVE; digit1<=NINE; digit2<=FIVE; digit3<=ONE; end
      16'd1596: begin digit0<=SIX; digit1<=NINE; digit2<=FIVE; digit3<=ONE; end
      16'd1597: begin digit0<=SEVEN; digit1<=NINE; digit2<=FIVE; digit3<=ONE; end
      16'd1598: begin digit0<=EIGHT; digit1<=NINE; digit2<=FIVE; digit3<=ONE; end
      16'd1599: begin digit0<=NINE; digit1<=NINE; digit2<=FIVE; digit3<=ONE; end
	  16'd1600: begin digit0<=ZERO; digit1<=ZERO; digit2<=SIX; digit3<=ONE; end
      16'd1601: begin digit0<=ONE; digit1<=ZERO; digit2<=SIX; digit3<=ONE; end
      16'd1602: begin digit0<=TWO; digit1<=ZERO; digit2<=SIX; digit3<=ONE; end
      16'd1603: begin digit0<=THREE; digit1<=ZERO; digit2<=SIX; digit3<=ONE; end
      16'd1604: begin digit0<=FOUR; digit1<=ZERO; digit2<=SIX; digit3<=ONE; end
      16'd1605: begin digit0<=FIVE; digit1<=ZERO; digit2<=SIX; digit3<=ONE; end
      16'd1606: begin digit0<=SIX; digit1<=ZERO; digit2<=SIX; digit3<=ONE; end
      16'd1607: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SIX; digit3<=ONE; end
      16'd1608: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SIX; digit3<=ONE; end
      16'd1609: begin digit0<=NINE; digit1<=ZERO; digit2<=SIX; digit3<=ONE; end
      16'd1610: begin digit0<=ZERO; digit1<=ONE; digit2<=SIX; digit3<=ONE; end
      16'd1611: begin digit0<=ONE; digit1<=ONE; digit2<=SIX; digit3<=ONE; end
      16'd1612: begin digit0<=TWO; digit1<=ONE; digit2<=SIX; digit3<=ONE; end
      16'd1613: begin digit0<=THREE; digit1<=ONE; digit2<=SIX; digit3<=ONE; end
      16'd1614: begin digit0<=FOUR; digit1<=ONE; digit2<=SIX; digit3<=ONE; end
      16'd1615: begin digit0<=FIVE; digit1<=ONE; digit2<=SIX; digit3<=ONE; end
      16'd1616: begin digit0<=SIX; digit1<=ONE; digit2<=SIX; digit3<=ONE; end
      16'd1617: begin digit0<=SEVEN; digit1<=ONE; digit2<=SIX; digit3<=ONE; end
      16'd1618: begin digit0<=EIGHT; digit1<=ONE; digit2<=SIX; digit3<=ONE; end
      16'd1619: begin digit0<=NINE; digit1<=ONE; digit2<=SIX; digit3<=ONE; end
      16'd1620: begin digit0<=ZERO; digit1<=TWO; digit2<=SIX; digit3<=ONE; end
      16'd1621: begin digit0<=ONE; digit1<=TWO; digit2<=SIX; digit3<=ONE; end
      16'd1622: begin digit0<=TWO; digit1<=TWO; digit2<=SIX; digit3<=ONE; end
      16'd1623: begin digit0<=THREE; digit1<=TWO; digit2<=SIX; digit3<=ONE; end
      16'd1624: begin digit0<=FOUR; digit1<=TWO; digit2<=SIX; digit3<=ONE; end
      16'd1625: begin digit0<=FIVE; digit1<=TWO; digit2<=SIX; digit3<=ONE; end
      16'd1626: begin digit0<=SIX; digit1<=TWO; digit2<=SIX; digit3<=ONE; end
      16'd1627: begin digit0<=SEVEN; digit1<=TWO; digit2<=SIX; digit3<=ONE; end
      16'd1628: begin digit0<=EIGHT; digit1<=TWO; digit2<=SIX; digit3<=ONE; end
      16'd1629: begin digit0<=NINE; digit1<=TWO; digit2<=SIX; digit3<=ONE; end
      16'd1630: begin digit0<=ZERO; digit1<=THREE; digit2<=SIX; digit3<=ONE; end
      16'd1631: begin digit0<=ONE; digit1<=THREE; digit2<=SIX; digit3<=ONE; end
      16'd1632: begin digit0<=TWO; digit1<=THREE; digit2<=SIX; digit3<=ONE; end
      16'd1633: begin digit0<=THREE; digit1<=THREE; digit2<=SIX; digit3<=ONE; end
      16'd1634: begin digit0<=FOUR; digit1<=THREE; digit2<=SIX; digit3<=ONE; end
      16'd1635: begin digit0<=FIVE; digit1<=THREE; digit2<=SIX; digit3<=ONE; end
      16'd1636: begin digit0<=SIX; digit1<=THREE; digit2<=SIX; digit3<=ONE; end
      16'd1637: begin digit0<=SEVEN; digit1<=THREE; digit2<=SIX; digit3<=ONE; end
      16'd1638: begin digit0<=EIGHT; digit1<=THREE; digit2<=SIX; digit3<=ONE; end
      16'd1639: begin digit0<=NINE; digit1<=THREE; digit2<=SIX; digit3<=ONE; end
      16'd1640: begin digit0<=ZERO; digit1<=FOUR; digit2<=SIX; digit3<=ONE; end
      16'd1641: begin digit0<=ONE; digit1<=FOUR; digit2<=SIX; digit3<=ONE; end
      16'd1642: begin digit0<=TWO; digit1<=FOUR; digit2<=SIX; digit3<=ONE; end
      16'd1643: begin digit0<=THREE; digit1<=FOUR; digit2<=SIX; digit3<=ONE; end
      16'd1644: begin digit0<=FOUR; digit1<=FOUR; digit2<=SIX; digit3<=ONE; end
      16'd1645: begin digit0<=FIVE; digit1<=FOUR; digit2<=SIX; digit3<=ONE; end
      16'd1646: begin digit0<=SIX; digit1<=FOUR; digit2<=SIX; digit3<=ONE; end
      16'd1647: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SIX; digit3<=ONE; end
      16'd1648: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SIX; digit3<=ONE; end
      16'd1649: begin digit0<=NINE; digit1<=FOUR; digit2<=SIX; digit3<=ONE; end
      16'd1650: begin digit0<=ZERO; digit1<=FIVE; digit2<=SIX; digit3<=ONE; end
      16'd1651: begin digit0<=ONE; digit1<=FIVE; digit2<=SIX; digit3<=ONE; end
      16'd1652: begin digit0<=TWO; digit1<=FIVE; digit2<=SIX; digit3<=ONE; end
      16'd1653: begin digit0<=THREE; digit1<=FIVE; digit2<=SIX; digit3<=ONE; end
      16'd1654: begin digit0<=FOUR; digit1<=FIVE; digit2<=SIX; digit3<=ONE; end
      16'd1655: begin digit0<=FIVE; digit1<=FIVE; digit2<=SIX; digit3<=ONE; end
      16'd1656: begin digit0<=SIX; digit1<=FIVE; digit2<=SIX; digit3<=ONE; end
      16'd1657: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SIX; digit3<=ONE; end
      16'd1658: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SIX; digit3<=ONE; end
      16'd1659: begin digit0<=NINE; digit1<=FIVE; digit2<=SIX; digit3<=ONE; end
      16'd1660: begin digit0<=ZERO; digit1<=SIX; digit2<=SIX; digit3<=ONE; end
      16'd1661: begin digit0<=ONE; digit1<=SIX; digit2<=SIX; digit3<=ONE; end
      16'd1662: begin digit0<=TWO; digit1<=SIX; digit2<=SIX; digit3<=ONE; end
      16'd1663: begin digit0<=THREE; digit1<=SIX; digit2<=SIX; digit3<=ONE; end
      16'd1664: begin digit0<=FOUR; digit1<=SIX; digit2<=SIX; digit3<=ONE; end
      16'd1665: begin digit0<=FIVE; digit1<=SIX; digit2<=SIX; digit3<=ONE; end
      16'd1666: begin digit0<=SIX; digit1<=SIX; digit2<=SIX; digit3<=ONE; end
      16'd1667: begin digit0<=SEVEN; digit1<=SIX; digit2<=SIX; digit3<=ONE; end
      16'd1668: begin digit0<=EIGHT; digit1<=SIX; digit2<=SIX; digit3<=ONE; end
      16'd1669: begin digit0<=NINE; digit1<=SIX; digit2<=SIX; digit3<=ONE; end
      16'd1670: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SIX; digit3<=ONE; end
      16'd1671: begin digit0<=ONE; digit1<=SEVEN; digit2<=SIX; digit3<=ONE; end
      16'd1672: begin digit0<=TWO; digit1<=SEVEN; digit2<=SIX; digit3<=ONE; end
      16'd1673: begin digit0<=THREE; digit1<=SEVEN; digit2<=SIX; digit3<=ONE; end
      16'd1674: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SIX; digit3<=ONE; end
      16'd1675: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SIX; digit3<=ONE; end
      16'd1676: begin digit0<=SIX; digit1<=SEVEN; digit2<=SIX; digit3<=ONE; end
      16'd1677: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SIX; digit3<=ONE; end
      16'd1678: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SIX; digit3<=ONE; end
      16'd1679: begin digit0<=NINE; digit1<=SEVEN; digit2<=SIX; digit3<=ONE; end
      16'd1680: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=ONE; end
      16'd1681: begin digit0<=ONE; digit1<=EIGHT; digit2<=SIX; digit3<=ONE; end
      16'd1682: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=ONE; end
      16'd1683: begin digit0<=THREE; digit1<=EIGHT; digit2<=SIX; digit3<=ONE; end
      16'd1684: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SIX; digit3<=ONE; end
      16'd1685: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SIX; digit3<=ONE; end
      16'd1686: begin digit0<=SIX; digit1<=EIGHT; digit2<=SIX; digit3<=ONE; end
      16'd1687: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SIX; digit3<=ONE; end
      16'd1688: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SIX; digit3<=ONE; end
      16'd1689: begin digit0<=NINE; digit1<=EIGHT; digit2<=SIX; digit3<=ONE; end
      16'd1690: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=ONE; end
      16'd1691: begin digit0<=ONE; digit1<=NINE; digit2<=SIX; digit3<=ONE; end
      16'd1692: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=ONE; end
      16'd1693: begin digit0<=THREE; digit1<=NINE; digit2<=SIX; digit3<=ONE; end
      16'd1694: begin digit0<=FOUR; digit1<=NINE; digit2<=SIX; digit3<=ONE; end
      16'd1695: begin digit0<=FIVE; digit1<=NINE; digit2<=SIX; digit3<=ONE; end
      16'd1696: begin digit0<=SIX; digit1<=NINE; digit2<=SIX; digit3<=ONE; end
      16'd1697: begin digit0<=SEVEN; digit1<=NINE; digit2<=SIX; digit3<=ONE; end
      16'd1698: begin digit0<=EIGHT; digit1<=NINE; digit2<=SIX; digit3<=ONE; end
      16'd1699: begin digit0<=NINE; digit1<=NINE; digit2<=SIX; digit3<=ONE; end
	  16'd1700: begin digit0<=ZERO; digit1<=ZERO; digit2<=SEVEN; digit3<=ONE; end
      16'd1701: begin digit0<=ONE; digit1<=ZERO; digit2<=SEVEN; digit3<=ONE; end
      16'd1702: begin digit0<=TWO; digit1<=ZERO; digit2<=SEVEN; digit3<=ONE; end
      16'd1703: begin digit0<=THREE; digit1<=ZERO; digit2<=SEVEN; digit3<=ONE; end
      16'd1704: begin digit0<=FOUR; digit1<=ZERO; digit2<=SEVEN; digit3<=ONE; end
      16'd1705: begin digit0<=FIVE; digit1<=ZERO; digit2<=SEVEN; digit3<=ONE; end
      16'd1706: begin digit0<=SIX; digit1<=ZERO; digit2<=SEVEN; digit3<=ONE; end
      16'd1707: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SEVEN; digit3<=ONE; end
      16'd1708: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SEVEN; digit3<=ONE; end
      16'd1709: begin digit0<=NINE; digit1<=ZERO; digit2<=SEVEN; digit3<=ONE; end
      16'd1710: begin digit0<=ZERO; digit1<=ONE; digit2<=SEVEN; digit3<=ONE; end
      16'd1711: begin digit0<=ONE; digit1<=ONE; digit2<=SEVEN; digit3<=ONE; end
      16'd1712: begin digit0<=TWO; digit1<=ONE; digit2<=SEVEN; digit3<=ONE; end
      16'd1713: begin digit0<=THREE; digit1<=ONE; digit2<=SEVEN; digit3<=ONE; end
      16'd1714: begin digit0<=FOUR; digit1<=ONE; digit2<=SEVEN; digit3<=ONE; end
      16'd1715: begin digit0<=FIVE; digit1<=ONE; digit2<=SEVEN; digit3<=ONE; end
      16'd1716: begin digit0<=SIX; digit1<=ONE; digit2<=SEVEN; digit3<=ONE; end
      16'd1717: begin digit0<=SEVEN; digit1<=ONE; digit2<=SEVEN; digit3<=ONE; end
      16'd1718: begin digit0<=EIGHT; digit1<=ONE; digit2<=SEVEN; digit3<=ONE; end
      16'd1719: begin digit0<=NINE; digit1<=ONE; digit2<=SEVEN; digit3<=ONE; end
      16'd1720: begin digit0<=ZERO; digit1<=TWO; digit2<=SEVEN; digit3<=ONE; end
      16'd1721: begin digit0<=ONE; digit1<=TWO; digit2<=SEVEN; digit3<=ONE; end
      16'd1722: begin digit0<=TWO; digit1<=TWO; digit2<=SEVEN; digit3<=ONE; end
      16'd1723: begin digit0<=THREE; digit1<=TWO; digit2<=SEVEN; digit3<=ONE; end
      16'd1724: begin digit0<=FOUR; digit1<=TWO; digit2<=SEVEN; digit3<=ONE; end
      16'd1725: begin digit0<=FIVE; digit1<=TWO; digit2<=SEVEN; digit3<=ONE; end
      16'd1726: begin digit0<=SIX; digit1<=TWO; digit2<=SEVEN; digit3<=ONE; end
      16'd1727: begin digit0<=SEVEN; digit1<=TWO; digit2<=SEVEN; digit3<=ONE; end
      16'd1728: begin digit0<=EIGHT; digit1<=TWO; digit2<=SEVEN; digit3<=ONE; end
      16'd1729: begin digit0<=NINE; digit1<=TWO; digit2<=SEVEN; digit3<=ONE; end
      16'd1730: begin digit0<=ZERO; digit1<=THREE; digit2<=SEVEN; digit3<=ONE; end
      16'd1731: begin digit0<=ONE; digit1<=THREE; digit2<=SEVEN; digit3<=ONE; end
      16'd1732: begin digit0<=TWO; digit1<=THREE; digit2<=SEVEN; digit3<=ONE; end
      16'd1733: begin digit0<=THREE; digit1<=THREE; digit2<=SEVEN; digit3<=ONE; end
      16'd1734: begin digit0<=FOUR; digit1<=THREE; digit2<=SEVEN; digit3<=ONE; end
      16'd1735: begin digit0<=FIVE; digit1<=THREE; digit2<=SEVEN; digit3<=ONE; end
      16'd1736: begin digit0<=SIX; digit1<=THREE; digit2<=SEVEN; digit3<=ONE; end
      16'd1737: begin digit0<=SEVEN; digit1<=THREE; digit2<=SEVEN; digit3<=ONE; end
      16'd1738: begin digit0<=EIGHT; digit1<=THREE; digit2<=SEVEN; digit3<=ONE; end
      16'd1739: begin digit0<=NINE; digit1<=THREE; digit2<=SEVEN; digit3<=ONE; end
      16'd1740: begin digit0<=ZERO; digit1<=FOUR; digit2<=SEVEN; digit3<=ONE; end
      16'd1741: begin digit0<=ONE; digit1<=FOUR; digit2<=SEVEN; digit3<=ONE; end
      16'd1742: begin digit0<=TWO; digit1<=FOUR; digit2<=SEVEN; digit3<=ONE; end
      16'd1743: begin digit0<=THREE; digit1<=FOUR; digit2<=SEVEN; digit3<=ONE; end
      16'd1744: begin digit0<=FOUR; digit1<=FOUR; digit2<=SEVEN; digit3<=ONE; end
      16'd1745: begin digit0<=FIVE; digit1<=FOUR; digit2<=SEVEN; digit3<=ONE; end
      16'd1746: begin digit0<=SIX; digit1<=FOUR; digit2<=SEVEN; digit3<=ONE; end
      16'd1747: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SEVEN; digit3<=ONE; end
      16'd1748: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SEVEN; digit3<=ONE; end
      16'd1749: begin digit0<=NINE; digit1<=FOUR; digit2<=SEVEN; digit3<=ONE; end
      16'd1750: begin digit0<=ZERO; digit1<=FIVE; digit2<=SEVEN; digit3<=ONE; end
      16'd1751: begin digit0<=ONE; digit1<=FIVE; digit2<=SEVEN; digit3<=ONE; end
      16'd1752: begin digit0<=TWO; digit1<=FIVE; digit2<=SEVEN; digit3<=ONE; end
      16'd1753: begin digit0<=THREE; digit1<=FIVE; digit2<=SEVEN; digit3<=ONE; end
      16'd1754: begin digit0<=FOUR; digit1<=FIVE; digit2<=SEVEN; digit3<=ONE; end
      16'd1755: begin digit0<=FIVE; digit1<=FIVE; digit2<=SEVEN; digit3<=ONE; end
      16'd1756: begin digit0<=SIX; digit1<=FIVE; digit2<=SEVEN; digit3<=ONE; end
      16'd1757: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SEVEN; digit3<=ONE; end
      16'd1758: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SEVEN; digit3<=ONE; end
      16'd1759: begin digit0<=NINE; digit1<=FIVE; digit2<=SEVEN; digit3<=ONE; end
      16'd1760: begin digit0<=ZERO; digit1<=SIX; digit2<=SEVEN; digit3<=ONE; end
      16'd1761: begin digit0<=ONE; digit1<=SIX; digit2<=SEVEN; digit3<=ONE; end
      16'd1762: begin digit0<=TWO; digit1<=SIX; digit2<=SEVEN; digit3<=ONE; end
      16'd1763: begin digit0<=THREE; digit1<=SIX; digit2<=SEVEN; digit3<=ONE; end
      16'd1764: begin digit0<=FOUR; digit1<=SIX; digit2<=SEVEN; digit3<=ONE; end
      16'd1765: begin digit0<=FIVE; digit1<=SIX; digit2<=SEVEN; digit3<=ONE; end
      16'd1766: begin digit0<=SIX; digit1<=SIX; digit2<=SEVEN; digit3<=ONE; end
      16'd1767: begin digit0<=SEVEN; digit1<=SIX; digit2<=SEVEN; digit3<=ONE; end
      16'd1768: begin digit0<=EIGHT; digit1<=SIX; digit2<=SEVEN; digit3<=ONE; end
      16'd1769: begin digit0<=NINE; digit1<=SIX; digit2<=SEVEN; digit3<=ONE; end
      16'd1770: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SEVEN; digit3<=ONE; end
      16'd1771: begin digit0<=ONE; digit1<=SEVEN; digit2<=SEVEN; digit3<=ONE; end
      16'd1772: begin digit0<=TWO; digit1<=SEVEN; digit2<=SEVEN; digit3<=ONE; end
      16'd1773: begin digit0<=THREE; digit1<=SEVEN; digit2<=SEVEN; digit3<=ONE; end
      16'd1774: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SEVEN; digit3<=ONE; end
      16'd1775: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SEVEN; digit3<=ONE; end
      16'd1776: begin digit0<=SIX; digit1<=SEVEN; digit2<=SEVEN; digit3<=ONE; end
      16'd1777: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SEVEN; digit3<=ONE; end
      16'd1778: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SEVEN; digit3<=ONE; end
      16'd1779: begin digit0<=NINE; digit1<=SEVEN; digit2<=SEVEN; digit3<=ONE; end
      16'd1780: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=ONE; end
      16'd1781: begin digit0<=ONE; digit1<=EIGHT; digit2<=SEVEN; digit3<=ONE; end
      16'd1782: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=ONE; end
      16'd1783: begin digit0<=THREE; digit1<=EIGHT; digit2<=SEVEN; digit3<=ONE; end
      16'd1784: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SEVEN; digit3<=ONE; end
      16'd1785: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SEVEN; digit3<=ONE; end
      16'd1786: begin digit0<=SIX; digit1<=EIGHT; digit2<=SEVEN; digit3<=ONE; end
      16'd1787: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SEVEN; digit3<=ONE; end
      16'd1788: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SEVEN; digit3<=ONE; end
      16'd1789: begin digit0<=NINE; digit1<=EIGHT; digit2<=SEVEN; digit3<=ONE; end
      16'd1790: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=ONE; end
      16'd1791: begin digit0<=ONE; digit1<=NINE; digit2<=SEVEN; digit3<=ONE; end
      16'd1792: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=ONE; end
      16'd1793: begin digit0<=THREE; digit1<=NINE; digit2<=SEVEN; digit3<=ONE; end
      16'd1794: begin digit0<=FOUR; digit1<=NINE; digit2<=SEVEN; digit3<=ONE; end
      16'd1795: begin digit0<=FIVE; digit1<=NINE; digit2<=SEVEN; digit3<=ONE; end
      16'd1796: begin digit0<=SIX; digit1<=NINE; digit2<=SEVEN; digit3<=ONE; end
      16'd1797: begin digit0<=SEVEN; digit1<=NINE; digit2<=SEVEN; digit3<=ONE; end
      16'd1798: begin digit0<=EIGHT; digit1<=NINE; digit2<=SEVEN; digit3<=ONE; end
      16'd1799: begin digit0<=NINE; digit1<=NINE; digit2<=SEVEN; digit3<=ONE; end
	  16'd1800: begin digit0<=ZERO; digit1<=ZERO; digit2<=EIGHT; digit3<=ONE; end
      16'd1801: begin digit0<=ONE; digit1<=ZERO; digit2<=EIGHT; digit3<=ONE; end
      16'd1802: begin digit0<=TWO; digit1<=ZERO; digit2<=EIGHT; digit3<=ONE; end
      16'd1803: begin digit0<=THREE; digit1<=ZERO; digit2<=EIGHT; digit3<=ONE; end
      16'd1804: begin digit0<=FOUR; digit1<=ZERO; digit2<=EIGHT; digit3<=ONE; end
      16'd1805: begin digit0<=FIVE; digit1<=ZERO; digit2<=EIGHT; digit3<=ONE; end
      16'd1806: begin digit0<=SIX; digit1<=ZERO; digit2<=EIGHT; digit3<=ONE; end
      16'd1807: begin digit0<=SEVEN; digit1<=ZERO; digit2<=EIGHT; digit3<=ONE; end
      16'd1808: begin digit0<=EIGHT; digit1<=ZERO; digit2<=EIGHT; digit3<=ONE; end
      16'd1809: begin digit0<=NINE; digit1<=ZERO; digit2<=EIGHT; digit3<=ONE; end
      16'd1810: begin digit0<=ZERO; digit1<=ONE; digit2<=EIGHT; digit3<=ONE; end
      16'd1811: begin digit0<=ONE; digit1<=ONE; digit2<=EIGHT; digit3<=ONE; end
      16'd1812: begin digit0<=TWO; digit1<=ONE; digit2<=EIGHT; digit3<=ONE; end
      16'd1813: begin digit0<=THREE; digit1<=ONE; digit2<=EIGHT; digit3<=ONE; end
      16'd1814: begin digit0<=FOUR; digit1<=ONE; digit2<=EIGHT; digit3<=ONE; end
      16'd1815: begin digit0<=FIVE; digit1<=ONE; digit2<=EIGHT; digit3<=ONE; end
      16'd1816: begin digit0<=SIX; digit1<=ONE; digit2<=EIGHT; digit3<=ONE; end
      16'd1817: begin digit0<=SEVEN; digit1<=ONE; digit2<=EIGHT; digit3<=ONE; end
      16'd1818: begin digit0<=EIGHT; digit1<=ONE; digit2<=EIGHT; digit3<=ONE; end
      16'd1819: begin digit0<=NINE; digit1<=ONE; digit2<=EIGHT; digit3<=ONE; end
      16'd1820: begin digit0<=ZERO; digit1<=TWO; digit2<=EIGHT; digit3<=ONE; end
      16'd1821: begin digit0<=ONE; digit1<=TWO; digit2<=EIGHT; digit3<=ONE; end
      16'd1822: begin digit0<=TWO; digit1<=TWO; digit2<=EIGHT; digit3<=ONE; end
      16'd1823: begin digit0<=THREE; digit1<=TWO; digit2<=EIGHT; digit3<=ONE; end
      16'd1824: begin digit0<=FOUR; digit1<=TWO; digit2<=EIGHT; digit3<=ONE; end
      16'd1825: begin digit0<=FIVE; digit1<=TWO; digit2<=EIGHT; digit3<=ONE; end
      16'd1826: begin digit0<=SIX; digit1<=TWO; digit2<=EIGHT; digit3<=ONE; end
      16'd1827: begin digit0<=SEVEN; digit1<=TWO; digit2<=EIGHT; digit3<=ONE; end
      16'd1828: begin digit0<=EIGHT; digit1<=TWO; digit2<=EIGHT; digit3<=ONE; end
      16'd1829: begin digit0<=NINE; digit1<=TWO; digit2<=EIGHT; digit3<=ONE; end
      16'd1830: begin digit0<=ZERO; digit1<=THREE; digit2<=EIGHT; digit3<=ONE; end
      16'd1831: begin digit0<=ONE; digit1<=THREE; digit2<=EIGHT; digit3<=ONE; end
      16'd1832: begin digit0<=TWO; digit1<=THREE; digit2<=EIGHT; digit3<=ONE; end
      16'd1833: begin digit0<=THREE; digit1<=THREE; digit2<=EIGHT; digit3<=ONE; end
      16'd1834: begin digit0<=FOUR; digit1<=THREE; digit2<=EIGHT; digit3<=ONE; end
      16'd1835: begin digit0<=FIVE; digit1<=THREE; digit2<=EIGHT; digit3<=ONE; end
      16'd1836: begin digit0<=SIX; digit1<=THREE; digit2<=EIGHT; digit3<=ONE; end
      16'd1837: begin digit0<=SEVEN; digit1<=THREE; digit2<=EIGHT; digit3<=ONE; end
      16'd1838: begin digit0<=EIGHT; digit1<=THREE; digit2<=EIGHT; digit3<=ONE; end
      16'd1839: begin digit0<=NINE; digit1<=THREE; digit2<=EIGHT; digit3<=ONE; end
      16'd1840: begin digit0<=ZERO; digit1<=FOUR; digit2<=EIGHT; digit3<=ONE; end
      16'd1841: begin digit0<=ONE; digit1<=FOUR; digit2<=EIGHT; digit3<=ONE; end
      16'd1842: begin digit0<=TWO; digit1<=FOUR; digit2<=EIGHT; digit3<=ONE; end
      16'd1843: begin digit0<=THREE; digit1<=FOUR; digit2<=EIGHT; digit3<=ONE; end
      16'd1844: begin digit0<=FOUR; digit1<=FOUR; digit2<=EIGHT; digit3<=ONE; end
      16'd1845: begin digit0<=FIVE; digit1<=FOUR; digit2<=EIGHT; digit3<=ONE; end
      16'd1846: begin digit0<=SIX; digit1<=FOUR; digit2<=EIGHT; digit3<=ONE; end
      16'd1847: begin digit0<=SEVEN; digit1<=FOUR; digit2<=EIGHT; digit3<=ONE; end
      16'd1848: begin digit0<=EIGHT; digit1<=FOUR; digit2<=EIGHT; digit3<=ONE; end
      16'd1849: begin digit0<=NINE; digit1<=FOUR; digit2<=EIGHT; digit3<=ONE; end
      16'd1850: begin digit0<=ZERO; digit1<=FIVE; digit2<=EIGHT; digit3<=ONE; end
      16'd1851: begin digit0<=ONE; digit1<=FIVE; digit2<=EIGHT; digit3<=ONE; end
      16'd1852: begin digit0<=TWO; digit1<=FIVE; digit2<=EIGHT; digit3<=ONE; end
      16'd1853: begin digit0<=THREE; digit1<=FIVE; digit2<=EIGHT; digit3<=ONE; end
      16'd1854: begin digit0<=FOUR; digit1<=FIVE; digit2<=EIGHT; digit3<=ONE; end
      16'd1855: begin digit0<=FIVE; digit1<=FIVE; digit2<=EIGHT; digit3<=ONE; end
      16'd1856: begin digit0<=SIX; digit1<=FIVE; digit2<=EIGHT; digit3<=ONE; end
      16'd1857: begin digit0<=SEVEN; digit1<=FIVE; digit2<=EIGHT; digit3<=ONE; end
      16'd1858: begin digit0<=EIGHT; digit1<=FIVE; digit2<=EIGHT; digit3<=ONE; end
      16'd1859: begin digit0<=NINE; digit1<=FIVE; digit2<=EIGHT; digit3<=ONE; end
      16'd1860: begin digit0<=ZERO; digit1<=SIX; digit2<=EIGHT; digit3<=ONE; end
      16'd1861: begin digit0<=ONE; digit1<=SIX; digit2<=EIGHT; digit3<=ONE; end
      16'd1862: begin digit0<=TWO; digit1<=SIX; digit2<=EIGHT; digit3<=ONE; end
      16'd1863: begin digit0<=THREE; digit1<=SIX; digit2<=EIGHT; digit3<=ONE; end
      16'd1864: begin digit0<=FOUR; digit1<=SIX; digit2<=EIGHT; digit3<=ONE; end
      16'd1865: begin digit0<=FIVE; digit1<=SIX; digit2<=EIGHT; digit3<=ONE; end
      16'd1866: begin digit0<=SIX; digit1<=SIX; digit2<=EIGHT; digit3<=ONE; end
      16'd1867: begin digit0<=SEVEN; digit1<=SIX; digit2<=EIGHT; digit3<=ONE; end
      16'd1868: begin digit0<=EIGHT; digit1<=SIX; digit2<=EIGHT; digit3<=ONE; end
      16'd1869: begin digit0<=NINE; digit1<=SIX; digit2<=EIGHT; digit3<=ONE; end
      16'd1870: begin digit0<=ZERO; digit1<=SEVEN; digit2<=EIGHT; digit3<=ONE; end
      16'd1871: begin digit0<=ONE; digit1<=SEVEN; digit2<=EIGHT; digit3<=ONE; end
      16'd1872: begin digit0<=TWO; digit1<=SEVEN; digit2<=EIGHT; digit3<=ONE; end
      16'd1873: begin digit0<=THREE; digit1<=SEVEN; digit2<=EIGHT; digit3<=ONE; end
      16'd1874: begin digit0<=FOUR; digit1<=SEVEN; digit2<=EIGHT; digit3<=ONE; end
      16'd1875: begin digit0<=FIVE; digit1<=SEVEN; digit2<=EIGHT; digit3<=ONE; end
      16'd1876: begin digit0<=SIX; digit1<=SEVEN; digit2<=EIGHT; digit3<=ONE; end
      16'd1877: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=EIGHT; digit3<=ONE; end
      16'd1878: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=EIGHT; digit3<=ONE; end
      16'd1879: begin digit0<=NINE; digit1<=SEVEN; digit2<=EIGHT; digit3<=ONE; end
      16'd1880: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=ONE; end
      16'd1881: begin digit0<=ONE; digit1<=EIGHT; digit2<=EIGHT; digit3<=ONE; end
      16'd1882: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=ONE; end
      16'd1883: begin digit0<=THREE; digit1<=EIGHT; digit2<=EIGHT; digit3<=ONE; end
      16'd1884: begin digit0<=FOUR; digit1<=EIGHT; digit2<=EIGHT; digit3<=ONE; end
      16'd1885: begin digit0<=FIVE; digit1<=EIGHT; digit2<=EIGHT; digit3<=ONE; end
      16'd1886: begin digit0<=SIX; digit1<=EIGHT; digit2<=EIGHT; digit3<=ONE; end
      16'd1887: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=EIGHT; digit3<=ONE; end
      16'd1888: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=EIGHT; digit3<=ONE; end
      16'd1889: begin digit0<=NINE; digit1<=EIGHT; digit2<=EIGHT; digit3<=ONE; end
      16'd1890: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=ONE; end
      16'd1891: begin digit0<=ONE; digit1<=NINE; digit2<=EIGHT; digit3<=ONE; end
      16'd1892: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=ONE; end
      16'd1893: begin digit0<=THREE; digit1<=NINE; digit2<=EIGHT; digit3<=ONE; end
      16'd1894: begin digit0<=FOUR; digit1<=NINE; digit2<=EIGHT; digit3<=ONE; end
      16'd1895: begin digit0<=FIVE; digit1<=NINE; digit2<=EIGHT; digit3<=ONE; end
      16'd1896: begin digit0<=SIX; digit1<=NINE; digit2<=EIGHT; digit3<=ONE; end
      16'd1897: begin digit0<=SEVEN; digit1<=NINE; digit2<=EIGHT; digit3<=ONE; end
      16'd1898: begin digit0<=EIGHT; digit1<=NINE; digit2<=EIGHT; digit3<=ONE; end
      16'd1899: begin digit0<=NINE; digit1<=NINE; digit2<=EIGHT; digit3<=ONE; end
	  16'd1900: begin digit0<=ZERO; digit1<=ZERO; digit2<=NINE; digit3<=ONE; end
      16'd1901: begin digit0<=ONE; digit1<=ZERO; digit2<=NINE; digit3<=ONE; end
      16'd1902: begin digit0<=TWO; digit1<=ZERO; digit2<=NINE; digit3<=ONE; end
      16'd1903: begin digit0<=THREE; digit1<=ZERO; digit2<=NINE; digit3<=ONE; end
      16'd1904: begin digit0<=FOUR; digit1<=ZERO; digit2<=NINE; digit3<=ONE; end
      16'd1905: begin digit0<=FIVE; digit1<=ZERO; digit2<=NINE; digit3<=ONE; end
      16'd1906: begin digit0<=SIX; digit1<=ZERO; digit2<=NINE; digit3<=ONE; end
      16'd1907: begin digit0<=SEVEN; digit1<=ZERO; digit2<=NINE; digit3<=ONE; end
      16'd1908: begin digit0<=EIGHT; digit1<=ZERO; digit2<=NINE; digit3<=ONE; end
      16'd1909: begin digit0<=NINE; digit1<=ZERO; digit2<=NINE; digit3<=ONE; end
      16'd1910: begin digit0<=ZERO; digit1<=ONE; digit2<=NINE; digit3<=ONE; end
      16'd1911: begin digit0<=ONE; digit1<=ONE; digit2<=NINE; digit3<=ONE; end
      16'd1912: begin digit0<=TWO; digit1<=ONE; digit2<=NINE; digit3<=ONE; end
      16'd1913: begin digit0<=THREE; digit1<=ONE; digit2<=NINE; digit3<=ONE; end
      16'd1914: begin digit0<=FOUR; digit1<=ONE; digit2<=NINE; digit3<=ONE; end
      16'd1915: begin digit0<=FIVE; digit1<=ONE; digit2<=NINE; digit3<=ONE; end
      16'd1916: begin digit0<=SIX; digit1<=ONE; digit2<=NINE; digit3<=ONE; end
      16'd1917: begin digit0<=SEVEN; digit1<=ONE; digit2<=NINE; digit3<=ONE; end
      16'd1918: begin digit0<=EIGHT; digit1<=ONE; digit2<=NINE; digit3<=ONE; end
      16'd1919: begin digit0<=NINE; digit1<=ONE; digit2<=NINE; digit3<=ONE; end
      16'd1920: begin digit0<=ZERO; digit1<=TWO; digit2<=NINE; digit3<=ONE; end
      16'd1921: begin digit0<=ONE; digit1<=TWO; digit2<=NINE; digit3<=ONE; end
      16'd1922: begin digit0<=TWO; digit1<=TWO; digit2<=NINE; digit3<=ONE; end
      16'd1923: begin digit0<=THREE; digit1<=TWO; digit2<=NINE; digit3<=ONE; end
      16'd1924: begin digit0<=FOUR; digit1<=TWO; digit2<=NINE; digit3<=ONE; end
      16'd1925: begin digit0<=FIVE; digit1<=TWO; digit2<=NINE; digit3<=ONE; end
      16'd1926: begin digit0<=SIX; digit1<=TWO; digit2<=NINE; digit3<=ONE; end
      16'd1927: begin digit0<=SEVEN; digit1<=TWO; digit2<=NINE; digit3<=ONE; end
      16'd1928: begin digit0<=EIGHT; digit1<=TWO; digit2<=NINE; digit3<=ONE; end
      16'd1929: begin digit0<=NINE; digit1<=TWO; digit2<=NINE; digit3<=ONE; end
      16'd1930: begin digit0<=ZERO; digit1<=THREE; digit2<=NINE; digit3<=ONE; end
      16'd1931: begin digit0<=ONE; digit1<=THREE; digit2<=NINE; digit3<=ONE; end
      16'd1932: begin digit0<=TWO; digit1<=THREE; digit2<=NINE; digit3<=ONE; end
      16'd1933: begin digit0<=THREE; digit1<=THREE; digit2<=NINE; digit3<=ONE; end
      16'd1934: begin digit0<=FOUR; digit1<=THREE; digit2<=NINE; digit3<=ONE; end
      16'd1935: begin digit0<=FIVE; digit1<=THREE; digit2<=NINE; digit3<=ONE; end
      16'd1936: begin digit0<=SIX; digit1<=THREE; digit2<=NINE; digit3<=ONE; end
      16'd1937: begin digit0<=SEVEN; digit1<=THREE; digit2<=NINE; digit3<=ONE; end
      16'd1938: begin digit0<=EIGHT; digit1<=THREE; digit2<=NINE; digit3<=ONE; end
      16'd1939: begin digit0<=NINE; digit1<=THREE; digit2<=NINE; digit3<=ONE; end
      16'd1940: begin digit0<=ZERO; digit1<=FOUR; digit2<=NINE; digit3<=ONE; end
      16'd1941: begin digit0<=ONE; digit1<=FOUR; digit2<=NINE; digit3<=ONE; end
      16'd1942: begin digit0<=TWO; digit1<=FOUR; digit2<=NINE; digit3<=ONE; end
      16'd1943: begin digit0<=THREE; digit1<=FOUR; digit2<=NINE; digit3<=ONE; end
      16'd1944: begin digit0<=FOUR; digit1<=FOUR; digit2<=NINE; digit3<=ONE; end
      16'd1945: begin digit0<=FIVE; digit1<=FOUR; digit2<=NINE; digit3<=ONE; end
      16'd1946: begin digit0<=SIX; digit1<=FOUR; digit2<=NINE; digit3<=ONE; end
      16'd1947: begin digit0<=SEVEN; digit1<=FOUR; digit2<=NINE; digit3<=ONE; end
      16'd1948: begin digit0<=EIGHT; digit1<=FOUR; digit2<=NINE; digit3<=ONE; end
      16'd1949: begin digit0<=NINE; digit1<=FOUR; digit2<=NINE; digit3<=ONE; end
      16'd1950: begin digit0<=ZERO; digit1<=FIVE; digit2<=NINE; digit3<=ONE; end
      16'd1951: begin digit0<=ONE; digit1<=FIVE; digit2<=NINE; digit3<=ONE; end
      16'd1952: begin digit0<=TWO; digit1<=FIVE; digit2<=NINE; digit3<=ONE; end
      16'd1953: begin digit0<=THREE; digit1<=FIVE; digit2<=NINE; digit3<=ONE; end
      16'd1954: begin digit0<=FOUR; digit1<=FIVE; digit2<=NINE; digit3<=ONE; end
      16'd1955: begin digit0<=FIVE; digit1<=FIVE; digit2<=NINE; digit3<=ONE; end
      16'd1956: begin digit0<=SIX; digit1<=FIVE; digit2<=NINE; digit3<=ONE; end
      16'd1957: begin digit0<=SEVEN; digit1<=FIVE; digit2<=NINE; digit3<=ONE; end
      16'd1958: begin digit0<=EIGHT; digit1<=FIVE; digit2<=NINE; digit3<=ONE; end
      16'd1959: begin digit0<=NINE; digit1<=FIVE; digit2<=NINE; digit3<=ONE; end
      16'd1960: begin digit0<=ZERO; digit1<=SIX; digit2<=NINE; digit3<=ONE; end
      16'd1961: begin digit0<=ONE; digit1<=SIX; digit2<=NINE; digit3<=ONE; end
      16'd1962: begin digit0<=TWO; digit1<=SIX; digit2<=NINE; digit3<=ONE; end
      16'd1963: begin digit0<=THREE; digit1<=SIX; digit2<=NINE; digit3<=ONE; end
      16'd1964: begin digit0<=FOUR; digit1<=SIX; digit2<=NINE; digit3<=ONE; end
      16'd1965: begin digit0<=FIVE; digit1<=SIX; digit2<=NINE; digit3<=ONE; end
      16'd1966: begin digit0<=SIX; digit1<=SIX; digit2<=NINE; digit3<=ONE; end
      16'd1967: begin digit0<=SEVEN; digit1<=SIX; digit2<=NINE; digit3<=ONE; end
      16'd1968: begin digit0<=EIGHT; digit1<=SIX; digit2<=NINE; digit3<=ONE; end
      16'd1969: begin digit0<=NINE; digit1<=SIX; digit2<=NINE; digit3<=ONE; end
      16'd1970: begin digit0<=ZERO; digit1<=SEVEN; digit2<=NINE; digit3<=ONE; end
      16'd1971: begin digit0<=ONE; digit1<=SEVEN; digit2<=NINE; digit3<=ONE; end
      16'd1972: begin digit0<=TWO; digit1<=SEVEN; digit2<=NINE; digit3<=ONE; end
      16'd1973: begin digit0<=THREE; digit1<=SEVEN; digit2<=NINE; digit3<=ONE; end
      16'd1974: begin digit0<=FOUR; digit1<=SEVEN; digit2<=NINE; digit3<=ONE; end
      16'd1975: begin digit0<=FIVE; digit1<=SEVEN; digit2<=NINE; digit3<=ONE; end
      16'd1976: begin digit0<=SIX; digit1<=SEVEN; digit2<=NINE; digit3<=ONE; end
      16'd1977: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=NINE; digit3<=ONE; end
      16'd1978: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=NINE; digit3<=ONE; end
      16'd1979: begin digit0<=NINE; digit1<=SEVEN; digit2<=NINE; digit3<=ONE; end
      16'd1980: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=ONE; end
      16'd1981: begin digit0<=ONE; digit1<=EIGHT; digit2<=NINE; digit3<=ONE; end
      16'd1982: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=ONE; end
      16'd1983: begin digit0<=THREE; digit1<=EIGHT; digit2<=NINE; digit3<=ONE; end
      16'd1984: begin digit0<=FOUR; digit1<=EIGHT; digit2<=NINE; digit3<=ONE; end
      16'd1985: begin digit0<=FIVE; digit1<=EIGHT; digit2<=NINE; digit3<=ONE; end
      16'd1986: begin digit0<=SIX; digit1<=EIGHT; digit2<=NINE; digit3<=ONE; end
      16'd1987: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=NINE; digit3<=ONE; end
      16'd1988: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=NINE; digit3<=ONE; end
      16'd1989: begin digit0<=NINE; digit1<=EIGHT; digit2<=NINE; digit3<=ONE; end
      16'd1990: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=ONE; end
      16'd1991: begin digit0<=ONE; digit1<=NINE; digit2<=NINE; digit3<=ONE; end
      16'd1992: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=ONE; end
      16'd1993: begin digit0<=THREE; digit1<=NINE; digit2<=NINE; digit3<=ONE; end
      16'd1994: begin digit0<=FOUR; digit1<=NINE; digit2<=NINE; digit3<=ONE; end
      16'd1995: begin digit0<=FIVE; digit1<=NINE; digit2<=NINE; digit3<=ONE; end
      16'd1996: begin digit0<=SIX; digit1<=NINE; digit2<=NINE; digit3<=ONE; end
      16'd1997: begin digit0<=SEVEN; digit1<=NINE; digit2<=NINE; digit3<=ONE; end
      16'd1998: begin digit0<=EIGHT; digit1<=NINE; digit2<=NINE; digit3<=ONE; end
      16'd1999: begin digit0<=NINE; digit1<=NINE; digit2<=NINE; digit3<=ONE; end
	  16'd2000: begin digit0<=ZERO; digit1<=ZERO; digit2<=ZERO; digit3<=TWO; end
      16'd2001: begin digit0<=ONE; digit1<=ZERO; digit2<=ZERO; digit3<=TWO; end
      16'd2002: begin digit0<=TWO; digit1<=ZERO; digit2<=ZERO; digit3<=TWO; end
      16'd2003: begin digit0<=THREE; digit1<=ZERO; digit2<=ZERO; digit3<=TWO; end
      16'd2004: begin digit0<=FOUR; digit1<=ZERO; digit2<=ZERO; digit3<=TWO; end
      16'd2005: begin digit0<=FIVE; digit1<=ZERO; digit2<=ZERO; digit3<=TWO; end
      16'd2006: begin digit0<=SIX; digit1<=ZERO; digit2<=ZERO; digit3<=TWO; end
      16'd2007: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ZERO; digit3<=TWO; end
      16'd2008: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ZERO; digit3<=TWO; end
      16'd2009: begin digit0<=NINE; digit1<=ZERO; digit2<=ZERO; digit3<=TWO; end
      16'd2010: begin digit0<=ZERO; digit1<=ONE; digit2<=ZERO; digit3<=TWO; end
      16'd2011: begin digit0<=ONE; digit1<=ONE; digit2<=ZERO; digit3<=TWO; end
      16'd2012: begin digit0<=TWO; digit1<=ONE; digit2<=ZERO; digit3<=TWO; end
      16'd2013: begin digit0<=THREE; digit1<=ONE; digit2<=ZERO; digit3<=TWO; end
      16'd2014: begin digit0<=FOUR; digit1<=ONE; digit2<=ZERO; digit3<=TWO; end
      16'd2015: begin digit0<=FIVE; digit1<=ONE; digit2<=ZERO; digit3<=TWO; end
      16'd2016: begin digit0<=SIX; digit1<=ONE; digit2<=ZERO; digit3<=TWO; end
      16'd2017: begin digit0<=SEVEN; digit1<=ONE; digit2<=ZERO; digit3<=TWO; end
      16'd2018: begin digit0<=EIGHT; digit1<=ONE; digit2<=ZERO; digit3<=TWO; end
      16'd2019: begin digit0<=NINE; digit1<=ONE; digit2<=ZERO; digit3<=TWO; end
      16'd2020: begin digit0<=ZERO; digit1<=TWO; digit2<=ZERO; digit3<=TWO; end
      16'd2021: begin digit0<=ONE; digit1<=TWO; digit2<=ZERO; digit3<=TWO; end
      16'd2022: begin digit0<=TWO; digit1<=TWO; digit2<=ZERO; digit3<=TWO; end
      16'd2023: begin digit0<=THREE; digit1<=TWO; digit2<=ZERO; digit3<=TWO; end
      16'd2024: begin digit0<=FOUR; digit1<=TWO; digit2<=ZERO; digit3<=TWO; end
      16'd2025: begin digit0<=FIVE; digit1<=TWO; digit2<=ZERO; digit3<=TWO; end
      16'd2026: begin digit0<=SIX; digit1<=TWO; digit2<=ZERO; digit3<=TWO; end
      16'd2027: begin digit0<=SEVEN; digit1<=TWO; digit2<=ZERO; digit3<=TWO; end
      16'd2028: begin digit0<=EIGHT; digit1<=TWO; digit2<=ZERO; digit3<=TWO; end
      16'd2029: begin digit0<=NINE; digit1<=TWO; digit2<=ZERO; digit3<=TWO; end
      16'd2030: begin digit0<=ZERO; digit1<=THREE; digit2<=ZERO; digit3<=TWO; end
      16'd2031: begin digit0<=ONE; digit1<=THREE; digit2<=ZERO; digit3<=TWO; end
      16'd2032: begin digit0<=TWO; digit1<=THREE; digit2<=ZERO; digit3<=TWO; end
      16'd2033: begin digit0<=THREE; digit1<=THREE; digit2<=ZERO; digit3<=TWO; end
      16'd2034: begin digit0<=FOUR; digit1<=THREE; digit2<=ZERO; digit3<=TWO; end
      16'd2035: begin digit0<=FIVE; digit1<=THREE; digit2<=ZERO; digit3<=TWO; end
      16'd2036: begin digit0<=SIX; digit1<=THREE; digit2<=ZERO; digit3<=TWO; end
      16'd2037: begin digit0<=SEVEN; digit1<=THREE; digit2<=ZERO; digit3<=TWO; end
      16'd2038: begin digit0<=EIGHT; digit1<=THREE; digit2<=ZERO; digit3<=TWO; end
      16'd2039: begin digit0<=NINE; digit1<=THREE; digit2<=ZERO; digit3<=TWO; end
      16'd2040: begin digit0<=ZERO; digit1<=FOUR; digit2<=ZERO; digit3<=TWO; end
      16'd2041: begin digit0<=ONE; digit1<=FOUR; digit2<=ZERO; digit3<=TWO; end
      16'd2042: begin digit0<=TWO; digit1<=FOUR; digit2<=ZERO; digit3<=TWO; end
      16'd2043: begin digit0<=THREE; digit1<=FOUR; digit2<=ZERO; digit3<=TWO; end
      16'd2044: begin digit0<=FOUR; digit1<=FOUR; digit2<=ZERO; digit3<=TWO; end
      16'd2045: begin digit0<=FIVE; digit1<=FOUR; digit2<=ZERO; digit3<=TWO; end
      16'd2046: begin digit0<=SIX; digit1<=FOUR; digit2<=ZERO; digit3<=TWO; end
      16'd2047: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ZERO; digit3<=TWO; end
      16'd2048: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ZERO; digit3<=TWO; end
      16'd2049: begin digit0<=NINE; digit1<=FOUR; digit2<=ZERO; digit3<=TWO; end
      16'd2050: begin digit0<=ZERO; digit1<=FIVE; digit2<=ZERO; digit3<=TWO; end
      16'd2051: begin digit0<=ONE; digit1<=FIVE; digit2<=ZERO; digit3<=TWO; end
      16'd2052: begin digit0<=TWO; digit1<=FIVE; digit2<=ZERO; digit3<=TWO; end
      16'd2053: begin digit0<=THREE; digit1<=FIVE; digit2<=ZERO; digit3<=TWO; end
      16'd2054: begin digit0<=FOUR; digit1<=FIVE; digit2<=ZERO; digit3<=TWO; end
      16'd2055: begin digit0<=FIVE; digit1<=FIVE; digit2<=ZERO; digit3<=TWO; end
      16'd2056: begin digit0<=SIX; digit1<=FIVE; digit2<=ZERO; digit3<=TWO; end
      16'd2057: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ZERO; digit3<=TWO; end
      16'd2058: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ZERO; digit3<=TWO; end
      16'd2059: begin digit0<=NINE; digit1<=FIVE; digit2<=ZERO; digit3<=TWO; end
      16'd2060: begin digit0<=ZERO; digit1<=SIX; digit2<=ZERO; digit3<=TWO; end
      16'd2061: begin digit0<=ONE; digit1<=SIX; digit2<=ZERO; digit3<=TWO; end
      16'd2062: begin digit0<=TWO; digit1<=SIX; digit2<=ZERO; digit3<=TWO; end
      16'd2063: begin digit0<=THREE; digit1<=SIX; digit2<=ZERO; digit3<=TWO; end
      16'd2064: begin digit0<=FOUR; digit1<=SIX; digit2<=ZERO; digit3<=TWO; end
      16'd2065: begin digit0<=FIVE; digit1<=SIX; digit2<=ZERO; digit3<=TWO; end
      16'd2066: begin digit0<=SIX; digit1<=SIX; digit2<=ZERO; digit3<=TWO; end
      16'd2067: begin digit0<=SEVEN; digit1<=SIX; digit2<=ZERO; digit3<=TWO; end
      16'd2068: begin digit0<=EIGHT; digit1<=SIX; digit2<=ZERO; digit3<=TWO; end
      16'd2069: begin digit0<=NINE; digit1<=SIX; digit2<=ZERO; digit3<=TWO; end
      16'd2070: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ZERO; digit3<=TWO; end
      16'd2071: begin digit0<=ONE; digit1<=SEVEN; digit2<=ZERO; digit3<=TWO; end
      16'd2072: begin digit0<=TWO; digit1<=SEVEN; digit2<=ZERO; digit3<=TWO; end
      16'd2073: begin digit0<=THREE; digit1<=SEVEN; digit2<=ZERO; digit3<=TWO; end
      16'd2074: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ZERO; digit3<=TWO; end
      16'd2075: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ZERO; digit3<=TWO; end
      16'd2076: begin digit0<=SIX; digit1<=SEVEN; digit2<=ZERO; digit3<=TWO; end
      16'd2077: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ZERO; digit3<=TWO; end
      16'd2078: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ZERO; digit3<=TWO; end
      16'd2079: begin digit0<=NINE; digit1<=SEVEN; digit2<=ZERO; digit3<=TWO; end
      16'd2080: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ZERO; digit3<=TWO; end
      16'd2081: begin digit0<=ONE; digit1<=EIGHT; digit2<=ZERO; digit3<=TWO; end
      16'd2082: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ZERO; digit3<=TWO; end
      16'd2083: begin digit0<=THREE; digit1<=EIGHT; digit2<=ZERO; digit3<=TWO; end
      16'd2084: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ZERO; digit3<=TWO; end
      16'd2085: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ZERO; digit3<=TWO; end
      16'd2086: begin digit0<=SIX; digit1<=EIGHT; digit2<=ZERO; digit3<=TWO; end
      16'd2087: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ZERO; digit3<=TWO; end
      16'd2088: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ZERO; digit3<=TWO; end
      16'd2089: begin digit0<=NINE; digit1<=EIGHT; digit2<=ZERO; digit3<=TWO; end
      16'd2090: begin digit0<=ZERO; digit1<=NINE; digit2<=ZERO; digit3<=TWO; end
      16'd2091: begin digit0<=ONE; digit1<=NINE; digit2<=ZERO; digit3<=TWO; end
      16'd2092: begin digit0<=ZERO; digit1<=NINE; digit2<=ZERO; digit3<=TWO; end
      16'd2093: begin digit0<=THREE; digit1<=NINE; digit2<=ZERO; digit3<=TWO; end
      16'd2094: begin digit0<=FOUR; digit1<=NINE; digit2<=ZERO; digit3<=TWO; end
      16'd2095: begin digit0<=FIVE; digit1<=NINE; digit2<=ZERO; digit3<=TWO; end
      16'd2096: begin digit0<=SIX; digit1<=NINE; digit2<=ZERO; digit3<=TWO; end
      16'd2097: begin digit0<=SEVEN; digit1<=NINE; digit2<=ZERO; digit3<=TWO; end
      16'd2098: begin digit0<=EIGHT; digit1<=NINE; digit2<=ZERO; digit3<=TWO; end
      16'd2099: begin digit0<=NINE; digit1<=NINE; digit2<=ZERO; digit3<=TWO; end
	  16'd2100: begin digit0<=ZERO; digit1<=ZERO; digit2<=ONE; digit3<=TWO; end
      16'd2101: begin digit0<=ONE; digit1<=ZERO; digit2<=ONE; digit3<=TWO; end
      16'd2102: begin digit0<=TWO; digit1<=ZERO; digit2<=ONE; digit3<=TWO; end
      16'd2103: begin digit0<=THREE; digit1<=ZERO; digit2<=ONE; digit3<=TWO; end
      16'd2104: begin digit0<=FOUR; digit1<=ZERO; digit2<=ONE; digit3<=TWO; end
      16'd2105: begin digit0<=FIVE; digit1<=ZERO; digit2<=ONE; digit3<=TWO; end
      16'd2106: begin digit0<=SIX; digit1<=ZERO; digit2<=ONE; digit3<=TWO; end
      16'd2107: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ONE; digit3<=TWO; end
      16'd2108: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ONE; digit3<=TWO; end
      16'd2109: begin digit0<=NINE; digit1<=ZERO; digit2<=ONE; digit3<=TWO; end
      16'd2110: begin digit0<=ZERO; digit1<=ONE; digit2<=ONE; digit3<=TWO; end
      16'd2111: begin digit0<=ONE; digit1<=ONE; digit2<=ONE; digit3<=TWO; end
      16'd2112: begin digit0<=TWO; digit1<=ONE; digit2<=ONE; digit3<=TWO; end
      16'd2113: begin digit0<=THREE; digit1<=ONE; digit2<=ONE; digit3<=TWO; end
      16'd2114: begin digit0<=FOUR; digit1<=ONE; digit2<=ONE; digit3<=TWO; end
      16'd2115: begin digit0<=FIVE; digit1<=ONE; digit2<=ONE; digit3<=TWO; end
      16'd2116: begin digit0<=SIX; digit1<=ONE; digit2<=ONE; digit3<=TWO; end
      16'd2117: begin digit0<=SEVEN; digit1<=ONE; digit2<=ONE; digit3<=TWO; end
      16'd2118: begin digit0<=EIGHT; digit1<=ONE; digit2<=ONE; digit3<=TWO; end
      16'd2119: begin digit0<=NINE; digit1<=ONE; digit2<=ONE; digit3<=TWO; end
      16'd2120: begin digit0<=ZERO; digit1<=TWO; digit2<=ONE; digit3<=TWO; end
      16'd2121: begin digit0<=ONE; digit1<=TWO; digit2<=ONE; digit3<=TWO; end
      16'd2122: begin digit0<=TWO; digit1<=TWO; digit2<=ONE; digit3<=TWO; end
      16'd2123: begin digit0<=THREE; digit1<=TWO; digit2<=ONE; digit3<=TWO; end
      16'd2124: begin digit0<=FOUR; digit1<=TWO; digit2<=ONE; digit3<=TWO; end
      16'd2125: begin digit0<=FIVE; digit1<=TWO; digit2<=ONE; digit3<=TWO; end
      16'd2126: begin digit0<=SIX; digit1<=TWO; digit2<=ONE; digit3<=TWO; end
      16'd2127: begin digit0<=SEVEN; digit1<=TWO; digit2<=ONE; digit3<=TWO; end
      16'd2128: begin digit0<=EIGHT; digit1<=TWO; digit2<=ONE; digit3<=TWO; end
      16'd2129: begin digit0<=NINE; digit1<=TWO; digit2<=ONE; digit3<=TWO; end
      16'd2130: begin digit0<=ZERO; digit1<=THREE; digit2<=ONE; digit3<=TWO; end
      16'd2131: begin digit0<=ONE; digit1<=THREE; digit2<=ONE; digit3<=TWO; end
      16'd2132: begin digit0<=TWO; digit1<=THREE; digit2<=ONE; digit3<=TWO; end
      16'd2133: begin digit0<=THREE; digit1<=THREE; digit2<=ONE; digit3<=TWO; end
      16'd2134: begin digit0<=FOUR; digit1<=THREE; digit2<=ONE; digit3<=TWO; end
      16'd2135: begin digit0<=FIVE; digit1<=THREE; digit2<=ONE; digit3<=TWO; end
      16'd2136: begin digit0<=SIX; digit1<=THREE; digit2<=ONE; digit3<=TWO; end
      16'd2137: begin digit0<=SEVEN; digit1<=THREE; digit2<=ONE; digit3<=TWO; end
      16'd2138: begin digit0<=EIGHT; digit1<=THREE; digit2<=ONE; digit3<=TWO; end
      16'd2139: begin digit0<=NINE; digit1<=THREE; digit2<=ONE; digit3<=TWO; end
      16'd2140: begin digit0<=ZERO; digit1<=FOUR; digit2<=ONE; digit3<=TWO; end
      16'd2141: begin digit0<=ONE; digit1<=FOUR; digit2<=ONE; digit3<=TWO; end
      16'd2142: begin digit0<=TWO; digit1<=FOUR; digit2<=ONE; digit3<=TWO; end
      16'd2143: begin digit0<=THREE; digit1<=FOUR; digit2<=ONE; digit3<=TWO; end
      16'd2144: begin digit0<=FOUR; digit1<=FOUR; digit2<=ONE; digit3<=TWO; end
      16'd2145: begin digit0<=FIVE; digit1<=FOUR; digit2<=ONE; digit3<=TWO; end
      16'd2146: begin digit0<=SIX; digit1<=FOUR; digit2<=ONE; digit3<=TWO; end
      16'd2147: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ONE; digit3<=TWO; end
      16'd2148: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ONE; digit3<=TWO; end
      16'd2149: begin digit0<=NINE; digit1<=FOUR; digit2<=ONE; digit3<=TWO; end
      16'd2150: begin digit0<=ZERO; digit1<=FIVE; digit2<=ONE; digit3<=TWO; end
      16'd2151: begin digit0<=ONE; digit1<=FIVE; digit2<=ONE; digit3<=TWO; end
      16'd2152: begin digit0<=TWO; digit1<=FIVE; digit2<=ONE; digit3<=TWO; end
      16'd2153: begin digit0<=THREE; digit1<=FIVE; digit2<=ONE; digit3<=TWO; end
      16'd2154: begin digit0<=FOUR; digit1<=FIVE; digit2<=ONE; digit3<=TWO; end
      16'd2155: begin digit0<=FIVE; digit1<=FIVE; digit2<=ONE; digit3<=TWO; end
      16'd2156: begin digit0<=SIX; digit1<=FIVE; digit2<=ONE; digit3<=TWO; end
      16'd2157: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ONE; digit3<=TWO; end
      16'd2158: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ONE; digit3<=TWO; end
      16'd2159: begin digit0<=NINE; digit1<=FIVE; digit2<=ONE; digit3<=TWO; end
      16'd2160: begin digit0<=ZERO; digit1<=SIX; digit2<=ONE; digit3<=TWO; end
      16'd2161: begin digit0<=ONE; digit1<=SIX; digit2<=ONE; digit3<=TWO; end
      16'd2162: begin digit0<=TWO; digit1<=SIX; digit2<=ONE; digit3<=TWO; end
      16'd2163: begin digit0<=THREE; digit1<=SIX; digit2<=ONE; digit3<=TWO; end
      16'd2164: begin digit0<=FOUR; digit1<=SIX; digit2<=ONE; digit3<=TWO; end
      16'd2165: begin digit0<=FIVE; digit1<=SIX; digit2<=ONE; digit3<=TWO; end
      16'd2166: begin digit0<=SIX; digit1<=SIX; digit2<=ONE; digit3<=TWO; end
      16'd2167: begin digit0<=SEVEN; digit1<=SIX; digit2<=ONE; digit3<=TWO; end
      16'd2168: begin digit0<=EIGHT; digit1<=SIX; digit2<=ONE; digit3<=TWO; end
      16'd2169: begin digit0<=NINE; digit1<=SIX; digit2<=ONE; digit3<=TWO; end
      16'd2170: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ONE; digit3<=TWO; end
      16'd2171: begin digit0<=ONE; digit1<=SEVEN; digit2<=ONE; digit3<=TWO; end
      16'd2172: begin digit0<=TWO; digit1<=SEVEN; digit2<=ONE; digit3<=TWO; end
      16'd2173: begin digit0<=THREE; digit1<=SEVEN; digit2<=ONE; digit3<=TWO; end
      16'd2174: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ONE; digit3<=TWO; end
      16'd2175: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ONE; digit3<=TWO; end
      16'd2176: begin digit0<=SIX; digit1<=SEVEN; digit2<=ONE; digit3<=TWO; end
      16'd2177: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ONE; digit3<=TWO; end
      16'd2178: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ONE; digit3<=TWO; end
      16'd2179: begin digit0<=NINE; digit1<=SEVEN; digit2<=ONE; digit3<=TWO; end
      16'd2180: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=TWO; end
      16'd2181: begin digit0<=ONE; digit1<=EIGHT; digit2<=ONE; digit3<=TWO; end
      16'd2182: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=TWO; end
      16'd2183: begin digit0<=THREE; digit1<=EIGHT; digit2<=ONE; digit3<=TWO; end
      16'd2184: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ONE; digit3<=TWO; end
      16'd2185: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ONE; digit3<=TWO; end
      16'd2186: begin digit0<=SIX; digit1<=EIGHT; digit2<=ONE; digit3<=TWO; end
      16'd2187: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ONE; digit3<=TWO; end
      16'd2188: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ONE; digit3<=TWO; end
      16'd2189: begin digit0<=NINE; digit1<=EIGHT; digit2<=ONE; digit3<=TWO; end
      16'd2190: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=TWO; end
      16'd2191: begin digit0<=ONE; digit1<=NINE; digit2<=ONE; digit3<=TWO; end
      16'd2192: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=TWO; end
      16'd2193: begin digit0<=THREE; digit1<=NINE; digit2<=ONE; digit3<=TWO; end
      16'd2194: begin digit0<=FOUR; digit1<=NINE; digit2<=ONE; digit3<=TWO; end
      16'd2195: begin digit0<=FIVE; digit1<=NINE; digit2<=ONE; digit3<=TWO; end
      16'd2196: begin digit0<=SIX; digit1<=NINE; digit2<=ONE; digit3<=TWO; end
      16'd2197: begin digit0<=SEVEN; digit1<=NINE; digit2<=ONE; digit3<=TWO; end
      16'd2198: begin digit0<=EIGHT; digit1<=NINE; digit2<=ONE; digit3<=TWO; end
      16'd2199: begin digit0<=NINE; digit1<=NINE; digit2<=ONE; digit3<=TWO; end
	  16'd2200: begin digit0<=ZERO; digit1<=ZERO; digit2<=TWO; digit3<=TWO; end
      16'd2201: begin digit0<=ONE; digit1<=ZERO; digit2<=TWO; digit3<=TWO; end
      16'd2202: begin digit0<=TWO; digit1<=ZERO; digit2<=TWO; digit3<=TWO; end
      16'd2203: begin digit0<=THREE; digit1<=ZERO; digit2<=TWO; digit3<=TWO; end
      16'd2204: begin digit0<=FOUR; digit1<=ZERO; digit2<=TWO; digit3<=TWO; end
      16'd2205: begin digit0<=FIVE; digit1<=ZERO; digit2<=TWO; digit3<=TWO; end
      16'd2206: begin digit0<=SIX; digit1<=ZERO; digit2<=TWO; digit3<=TWO; end
      16'd2207: begin digit0<=SEVEN; digit1<=ZERO; digit2<=TWO; digit3<=TWO; end
      16'd2208: begin digit0<=EIGHT; digit1<=ZERO; digit2<=TWO; digit3<=TWO; end
      16'd2209: begin digit0<=NINE; digit1<=ZERO; digit2<=TWO; digit3<=TWO; end
      16'd2210: begin digit0<=ZERO; digit1<=ONE; digit2<=TWO; digit3<=TWO; end
      16'd2211: begin digit0<=ONE; digit1<=ONE; digit2<=TWO; digit3<=TWO; end
      16'd2212: begin digit0<=TWO; digit1<=ONE; digit2<=TWO; digit3<=TWO; end
      16'd2213: begin digit0<=THREE; digit1<=ONE; digit2<=TWO; digit3<=TWO; end
      16'd2214: begin digit0<=FOUR; digit1<=ONE; digit2<=TWO; digit3<=TWO; end
      16'd2215: begin digit0<=FIVE; digit1<=ONE; digit2<=TWO; digit3<=TWO; end
      16'd2216: begin digit0<=SIX; digit1<=ONE; digit2<=TWO; digit3<=TWO; end
      16'd2217: begin digit0<=SEVEN; digit1<=ONE; digit2<=TWO; digit3<=TWO; end
      16'd2218: begin digit0<=EIGHT; digit1<=ONE; digit2<=TWO; digit3<=TWO; end
      16'd2219: begin digit0<=NINE; digit1<=ONE; digit2<=TWO; digit3<=TWO; end
      16'd2220: begin digit0<=ZERO; digit1<=TWO; digit2<=TWO; digit3<=TWO; end
      16'd2221: begin digit0<=ONE; digit1<=TWO; digit2<=TWO; digit3<=TWO; end
      16'd2222: begin digit0<=TWO; digit1<=TWO; digit2<=TWO; digit3<=TWO; end
      16'd2223: begin digit0<=THREE; digit1<=TWO; digit2<=TWO; digit3<=TWO; end
      16'd2224: begin digit0<=FOUR; digit1<=TWO; digit2<=TWO; digit3<=TWO; end
      16'd2225: begin digit0<=FIVE; digit1<=TWO; digit2<=TWO; digit3<=TWO; end
      16'd2226: begin digit0<=SIX; digit1<=TWO; digit2<=TWO; digit3<=TWO; end
      16'd2227: begin digit0<=SEVEN; digit1<=TWO; digit2<=TWO; digit3<=TWO; end
      16'd2228: begin digit0<=EIGHT; digit1<=TWO; digit2<=TWO; digit3<=TWO; end
      16'd2229: begin digit0<=NINE; digit1<=TWO; digit2<=TWO; digit3<=TWO; end
      16'd2230: begin digit0<=ZERO; digit1<=THREE; digit2<=TWO; digit3<=TWO; end
      16'd2231: begin digit0<=ONE; digit1<=THREE; digit2<=TWO; digit3<=TWO; end
      16'd2232: begin digit0<=TWO; digit1<=THREE; digit2<=TWO; digit3<=TWO; end
      16'd2233: begin digit0<=THREE; digit1<=THREE; digit2<=TWO; digit3<=TWO; end
      16'd2234: begin digit0<=FOUR; digit1<=THREE; digit2<=TWO; digit3<=TWO; end
      16'd2235: begin digit0<=FIVE; digit1<=THREE; digit2<=TWO; digit3<=TWO; end
      16'd2236: begin digit0<=SIX; digit1<=THREE; digit2<=TWO; digit3<=TWO; end
      16'd2237: begin digit0<=SEVEN; digit1<=THREE; digit2<=TWO; digit3<=TWO; end
      16'd2238: begin digit0<=EIGHT; digit1<=THREE; digit2<=TWO; digit3<=TWO; end
      16'd2239: begin digit0<=NINE; digit1<=THREE; digit2<=TWO; digit3<=TWO; end
      16'd2240: begin digit0<=ZERO; digit1<=FOUR; digit2<=TWO; digit3<=TWO; end
      16'd2241: begin digit0<=ONE; digit1<=FOUR; digit2<=TWO; digit3<=TWO; end
      16'd2242: begin digit0<=TWO; digit1<=FOUR; digit2<=TWO; digit3<=TWO; end
      16'd2243: begin digit0<=THREE; digit1<=FOUR; digit2<=TWO; digit3<=TWO; end
      16'd2244: begin digit0<=FOUR; digit1<=FOUR; digit2<=TWO; digit3<=TWO; end
      16'd2245: begin digit0<=FIVE; digit1<=FOUR; digit2<=TWO; digit3<=TWO; end
      16'd2246: begin digit0<=SIX; digit1<=FOUR; digit2<=TWO; digit3<=TWO; end
      16'd2247: begin digit0<=SEVEN; digit1<=FOUR; digit2<=TWO; digit3<=TWO; end
      16'd2248: begin digit0<=EIGHT; digit1<=FOUR; digit2<=TWO; digit3<=TWO; end
      16'd2249: begin digit0<=NINE; digit1<=FOUR; digit2<=TWO; digit3<=TWO; end
      16'd2250: begin digit0<=ZERO; digit1<=FIVE; digit2<=TWO; digit3<=TWO; end
      16'd2251: begin digit0<=ONE; digit1<=FIVE; digit2<=TWO; digit3<=TWO; end
      16'd2252: begin digit0<=TWO; digit1<=FIVE; digit2<=TWO; digit3<=TWO; end
      16'd2253: begin digit0<=THREE; digit1<=FIVE; digit2<=TWO; digit3<=TWO; end
      16'd2254: begin digit0<=FOUR; digit1<=FIVE; digit2<=TWO; digit3<=TWO; end
      16'd2255: begin digit0<=FIVE; digit1<=FIVE; digit2<=TWO; digit3<=TWO; end
      16'd2256: begin digit0<=SIX; digit1<=FIVE; digit2<=TWO; digit3<=TWO; end
      16'd2257: begin digit0<=SEVEN; digit1<=FIVE; digit2<=TWO; digit3<=TWO; end
      16'd2258: begin digit0<=EIGHT; digit1<=FIVE; digit2<=TWO; digit3<=TWO; end
      16'd2259: begin digit0<=NINE; digit1<=FIVE; digit2<=TWO; digit3<=TWO; end
      16'd2260: begin digit0<=ZERO; digit1<=SIX; digit2<=TWO; digit3<=TWO; end
      16'd2261: begin digit0<=ONE; digit1<=SIX; digit2<=TWO; digit3<=TWO; end
      16'd2262: begin digit0<=TWO; digit1<=SIX; digit2<=TWO; digit3<=TWO; end
      16'd2263: begin digit0<=THREE; digit1<=SIX; digit2<=TWO; digit3<=TWO; end
      16'd2264: begin digit0<=FOUR; digit1<=SIX; digit2<=TWO; digit3<=TWO; end
      16'd2265: begin digit0<=FIVE; digit1<=SIX; digit2<=TWO; digit3<=TWO; end
      16'd2266: begin digit0<=SIX; digit1<=SIX; digit2<=TWO; digit3<=TWO; end
      16'd2267: begin digit0<=SEVEN; digit1<=SIX; digit2<=TWO; digit3<=TWO; end
      16'd2268: begin digit0<=EIGHT; digit1<=SIX; digit2<=TWO; digit3<=TWO; end
      16'd2269: begin digit0<=NINE; digit1<=SIX; digit2<=TWO; digit3<=TWO; end
      16'd2270: begin digit0<=ZERO; digit1<=SEVEN; digit2<=TWO; digit3<=TWO; end
      16'd2271: begin digit0<=ONE; digit1<=SEVEN; digit2<=TWO; digit3<=TWO; end
      16'd2272: begin digit0<=TWO; digit1<=SEVEN; digit2<=TWO; digit3<=TWO; end
      16'd2273: begin digit0<=THREE; digit1<=SEVEN; digit2<=TWO; digit3<=TWO; end
      16'd2274: begin digit0<=FOUR; digit1<=SEVEN; digit2<=TWO; digit3<=TWO; end
      16'd2275: begin digit0<=FIVE; digit1<=SEVEN; digit2<=TWO; digit3<=TWO; end
      16'd2276: begin digit0<=SIX; digit1<=SEVEN; digit2<=TWO; digit3<=TWO; end
      16'd2277: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=TWO; digit3<=TWO; end
      16'd2278: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=TWO; digit3<=TWO; end
      16'd2279: begin digit0<=NINE; digit1<=SEVEN; digit2<=TWO; digit3<=TWO; end
      16'd2280: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=TWO; end
      16'd2281: begin digit0<=ONE; digit1<=EIGHT; digit2<=TWO; digit3<=TWO; end
      16'd2282: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=TWO; end
      16'd2283: begin digit0<=THREE; digit1<=EIGHT; digit2<=TWO; digit3<=TWO; end
      16'd2284: begin digit0<=FOUR; digit1<=EIGHT; digit2<=TWO; digit3<=TWO; end
      16'd2285: begin digit0<=FIVE; digit1<=EIGHT; digit2<=TWO; digit3<=TWO; end
      16'd2286: begin digit0<=SIX; digit1<=EIGHT; digit2<=TWO; digit3<=TWO; end
      16'd2287: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=TWO; digit3<=TWO; end
      16'd2288: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=TWO; digit3<=TWO; end
      16'd2289: begin digit0<=NINE; digit1<=EIGHT; digit2<=TWO; digit3<=TWO; end
      16'd2290: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=TWO; end
      16'd2291: begin digit0<=ONE; digit1<=NINE; digit2<=TWO; digit3<=TWO; end
      16'd2292: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=TWO; end
      16'd2293: begin digit0<=THREE; digit1<=NINE; digit2<=TWO; digit3<=TWO; end
      16'd2294: begin digit0<=FOUR; digit1<=NINE; digit2<=TWO; digit3<=TWO; end
      16'd2295: begin digit0<=FIVE; digit1<=NINE; digit2<=TWO; digit3<=TWO; end
      16'd2296: begin digit0<=SIX; digit1<=NINE; digit2<=TWO; digit3<=TWO; end
      16'd2297: begin digit0<=SEVEN; digit1<=NINE; digit2<=TWO; digit3<=TWO; end
      16'd2298: begin digit0<=EIGHT; digit1<=NINE; digit2<=TWO; digit3<=TWO; end
      16'd2299: begin digit0<=NINE; digit1<=NINE; digit2<=TWO; digit3<=TWO; end
	  16'd2300: begin digit0<=ZERO; digit1<=ZERO; digit2<=THREE; digit3<=TWO; end
      16'd2301: begin digit0<=ONE; digit1<=ZERO; digit2<=THREE; digit3<=TWO; end
      16'd2302: begin digit0<=TWO; digit1<=ZERO; digit2<=THREE; digit3<=TWO; end
      16'd2303: begin digit0<=THREE; digit1<=ZERO; digit2<=THREE; digit3<=TWO; end
      16'd2304: begin digit0<=FOUR; digit1<=ZERO; digit2<=THREE; digit3<=TWO; end
      16'd2305: begin digit0<=FIVE; digit1<=ZERO; digit2<=THREE; digit3<=TWO; end
      16'd2306: begin digit0<=SIX; digit1<=ZERO; digit2<=THREE; digit3<=TWO; end
      16'd2307: begin digit0<=SEVEN; digit1<=ZERO; digit2<=THREE; digit3<=TWO; end
      16'd2308: begin digit0<=EIGHT; digit1<=ZERO; digit2<=THREE; digit3<=TWO; end
      16'd2309: begin digit0<=NINE; digit1<=ZERO; digit2<=THREE; digit3<=TWO; end
      16'd2310: begin digit0<=ZERO; digit1<=ONE; digit2<=THREE; digit3<=TWO; end
      16'd2311: begin digit0<=ONE; digit1<=ONE; digit2<=THREE; digit3<=TWO; end
      16'd2312: begin digit0<=TWO; digit1<=ONE; digit2<=THREE; digit3<=TWO; end
      16'd2313: begin digit0<=THREE; digit1<=ONE; digit2<=THREE; digit3<=TWO; end
      16'd2314: begin digit0<=FOUR; digit1<=ONE; digit2<=THREE; digit3<=TWO; end
      16'd2315: begin digit0<=FIVE; digit1<=ONE; digit2<=THREE; digit3<=TWO; end
      16'd2316: begin digit0<=SIX; digit1<=ONE; digit2<=THREE; digit3<=TWO; end
      16'd2317: begin digit0<=SEVEN; digit1<=ONE; digit2<=THREE; digit3<=TWO; end
      16'd2318: begin digit0<=EIGHT; digit1<=ONE; digit2<=THREE; digit3<=TWO; end
      16'd2319: begin digit0<=NINE; digit1<=ONE; digit2<=THREE; digit3<=TWO; end
      16'd2320: begin digit0<=ZERO; digit1<=TWO; digit2<=THREE; digit3<=TWO; end
      16'd2321: begin digit0<=ONE; digit1<=TWO; digit2<=THREE; digit3<=TWO; end
      16'd2322: begin digit0<=TWO; digit1<=TWO; digit2<=THREE; digit3<=TWO; end
      16'd2323: begin digit0<=THREE; digit1<=TWO; digit2<=THREE; digit3<=TWO; end
      16'd2324: begin digit0<=FOUR; digit1<=TWO; digit2<=THREE; digit3<=TWO; end
      16'd2325: begin digit0<=FIVE; digit1<=TWO; digit2<=THREE; digit3<=TWO; end
      16'd2326: begin digit0<=SIX; digit1<=TWO; digit2<=THREE; digit3<=TWO; end
      16'd2327: begin digit0<=SEVEN; digit1<=TWO; digit2<=THREE; digit3<=TWO; end
      16'd2328: begin digit0<=EIGHT; digit1<=TWO; digit2<=THREE; digit3<=TWO; end
      16'd2329: begin digit0<=NINE; digit1<=TWO; digit2<=THREE; digit3<=TWO; end
      16'd2330: begin digit0<=ZERO; digit1<=THREE; digit2<=THREE; digit3<=TWO; end
      16'd2331: begin digit0<=ONE; digit1<=THREE; digit2<=THREE; digit3<=TWO; end
      16'd2332: begin digit0<=TWO; digit1<=THREE; digit2<=THREE; digit3<=TWO; end
      16'd2333: begin digit0<=THREE; digit1<=THREE; digit2<=THREE; digit3<=TWO; end
      16'd2334: begin digit0<=FOUR; digit1<=THREE; digit2<=THREE; digit3<=TWO; end
      16'd2335: begin digit0<=FIVE; digit1<=THREE; digit2<=THREE; digit3<=TWO; end
      16'd2336: begin digit0<=SIX; digit1<=THREE; digit2<=THREE; digit3<=TWO; end
      16'd2337: begin digit0<=SEVEN; digit1<=THREE; digit2<=THREE; digit3<=TWO; end
      16'd2338: begin digit0<=EIGHT; digit1<=THREE; digit2<=THREE; digit3<=TWO; end
      16'd2339: begin digit0<=NINE; digit1<=THREE; digit2<=THREE; digit3<=TWO; end
      16'd2340: begin digit0<=ZERO; digit1<=FOUR; digit2<=THREE; digit3<=TWO; end
      16'd2341: begin digit0<=ONE; digit1<=FOUR; digit2<=THREE; digit3<=TWO; end
      16'd2342: begin digit0<=TWO; digit1<=FOUR; digit2<=THREE; digit3<=TWO; end
      16'd2343: begin digit0<=THREE; digit1<=FOUR; digit2<=THREE; digit3<=TWO; end
      16'd2344: begin digit0<=FOUR; digit1<=FOUR; digit2<=THREE; digit3<=TWO; end
      16'd2345: begin digit0<=FIVE; digit1<=FOUR; digit2<=THREE; digit3<=TWO; end
      16'd2346: begin digit0<=SIX; digit1<=FOUR; digit2<=THREE; digit3<=TWO; end
      16'd2347: begin digit0<=SEVEN; digit1<=FOUR; digit2<=THREE; digit3<=TWO; end
      16'd2348: begin digit0<=EIGHT; digit1<=FOUR; digit2<=THREE; digit3<=TWO; end
      16'd2349: begin digit0<=NINE; digit1<=FOUR; digit2<=THREE; digit3<=TWO; end
      16'd2350: begin digit0<=ZERO; digit1<=FIVE; digit2<=THREE; digit3<=TWO; end
      16'd2351: begin digit0<=ONE; digit1<=FIVE; digit2<=THREE; digit3<=TWO; end
      16'd2352: begin digit0<=TWO; digit1<=FIVE; digit2<=THREE; digit3<=TWO; end
      16'd2353: begin digit0<=THREE; digit1<=FIVE; digit2<=THREE; digit3<=TWO; end
      16'd2354: begin digit0<=FOUR; digit1<=FIVE; digit2<=THREE; digit3<=TWO; end
      16'd2355: begin digit0<=FIVE; digit1<=FIVE; digit2<=THREE; digit3<=TWO; end
      16'd2356: begin digit0<=SIX; digit1<=FIVE; digit2<=THREE; digit3<=TWO; end
      16'd2357: begin digit0<=SEVEN; digit1<=FIVE; digit2<=THREE; digit3<=TWO; end
      16'd2358: begin digit0<=EIGHT; digit1<=FIVE; digit2<=THREE; digit3<=TWO; end
      16'd2359: begin digit0<=NINE; digit1<=FIVE; digit2<=THREE; digit3<=TWO; end
      16'd2360: begin digit0<=ZERO; digit1<=SIX; digit2<=THREE; digit3<=TWO; end
      16'd2361: begin digit0<=ONE; digit1<=SIX; digit2<=THREE; digit3<=TWO; end
      16'd2362: begin digit0<=TWO; digit1<=SIX; digit2<=THREE; digit3<=TWO; end
      16'd2363: begin digit0<=THREE; digit1<=SIX; digit2<=THREE; digit3<=TWO; end
      16'd2364: begin digit0<=FOUR; digit1<=SIX; digit2<=THREE; digit3<=TWO; end
      16'd2365: begin digit0<=FIVE; digit1<=SIX; digit2<=THREE; digit3<=TWO; end
      16'd2366: begin digit0<=SIX; digit1<=SIX; digit2<=THREE; digit3<=TWO; end
      16'd2367: begin digit0<=SEVEN; digit1<=SIX; digit2<=THREE; digit3<=TWO; end
      16'd2368: begin digit0<=EIGHT; digit1<=SIX; digit2<=THREE; digit3<=TWO; end
      16'd2369: begin digit0<=NINE; digit1<=SIX; digit2<=THREE; digit3<=TWO; end
      16'd2370: begin digit0<=ZERO; digit1<=SEVEN; digit2<=THREE; digit3<=TWO; end
      16'd2371: begin digit0<=ONE; digit1<=SEVEN; digit2<=THREE; digit3<=TWO; end
      16'd2372: begin digit0<=TWO; digit1<=SEVEN; digit2<=THREE; digit3<=TWO; end
      16'd2373: begin digit0<=THREE; digit1<=SEVEN; digit2<=THREE; digit3<=TWO; end
      16'd2374: begin digit0<=FOUR; digit1<=SEVEN; digit2<=THREE; digit3<=TWO; end
      16'd2375: begin digit0<=FIVE; digit1<=SEVEN; digit2<=THREE; digit3<=TWO; end
      16'd2376: begin digit0<=SIX; digit1<=SEVEN; digit2<=THREE; digit3<=TWO; end
      16'd2377: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=THREE; digit3<=TWO; end
      16'd2378: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=THREE; digit3<=TWO; end
      16'd2379: begin digit0<=NINE; digit1<=SEVEN; digit2<=THREE; digit3<=TWO; end
      16'd2380: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=TWO; end
      16'd2381: begin digit0<=ONE; digit1<=EIGHT; digit2<=THREE; digit3<=TWO; end
      16'd2382: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=TWO; end
      16'd2383: begin digit0<=THREE; digit1<=EIGHT; digit2<=THREE; digit3<=TWO; end
      16'd2384: begin digit0<=FOUR; digit1<=EIGHT; digit2<=THREE; digit3<=TWO; end
      16'd2385: begin digit0<=FIVE; digit1<=EIGHT; digit2<=THREE; digit3<=TWO; end
      16'd2386: begin digit0<=SIX; digit1<=EIGHT; digit2<=THREE; digit3<=TWO; end
      16'd2387: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=THREE; digit3<=TWO; end
      16'd2388: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=THREE; digit3<=TWO; end
      16'd2389: begin digit0<=NINE; digit1<=EIGHT; digit2<=THREE; digit3<=TWO; end
      16'd2390: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=TWO; end
      16'd2391: begin digit0<=ONE; digit1<=NINE; digit2<=THREE; digit3<=TWO; end
      16'd2392: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=TWO; end
      16'd2393: begin digit0<=THREE; digit1<=NINE; digit2<=THREE; digit3<=TWO; end
      16'd2394: begin digit0<=FOUR; digit1<=NINE; digit2<=THREE; digit3<=TWO; end
      16'd2395: begin digit0<=FIVE; digit1<=NINE; digit2<=THREE; digit3<=TWO; end
      16'd2396: begin digit0<=SIX; digit1<=NINE; digit2<=THREE; digit3<=TWO; end
      16'd2397: begin digit0<=SEVEN; digit1<=NINE; digit2<=THREE; digit3<=TWO; end
      16'd2398: begin digit0<=EIGHT; digit1<=NINE; digit2<=THREE; digit3<=TWO; end
      16'd2399: begin digit0<=NINE; digit1<=NINE; digit2<=THREE; digit3<=TWO; end
	  16'd2400: begin digit0<=ZERO; digit1<=ZERO; digit2<=FOUR; digit3<=TWO; end
      16'd2401: begin digit0<=ONE; digit1<=ZERO; digit2<=FOUR; digit3<=TWO; end
      16'd2402: begin digit0<=TWO; digit1<=ZERO; digit2<=FOUR; digit3<=TWO; end
      16'd2403: begin digit0<=THREE; digit1<=ZERO; digit2<=FOUR; digit3<=TWO; end
      16'd2404: begin digit0<=FOUR; digit1<=ZERO; digit2<=FOUR; digit3<=TWO; end
      16'd2405: begin digit0<=FIVE; digit1<=ZERO; digit2<=FOUR; digit3<=TWO; end
      16'd2406: begin digit0<=SIX; digit1<=ZERO; digit2<=FOUR; digit3<=TWO; end
      16'd2407: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FOUR; digit3<=TWO; end
      16'd2408: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FOUR; digit3<=TWO; end
      16'd2409: begin digit0<=NINE; digit1<=ZERO; digit2<=FOUR; digit3<=TWO; end
      16'd2410: begin digit0<=ZERO; digit1<=ONE; digit2<=FOUR; digit3<=TWO; end
      16'd2411: begin digit0<=ONE; digit1<=ONE; digit2<=FOUR; digit3<=TWO; end
      16'd2412: begin digit0<=TWO; digit1<=ONE; digit2<=FOUR; digit3<=TWO; end
      16'd2413: begin digit0<=THREE; digit1<=ONE; digit2<=FOUR; digit3<=TWO; end
      16'd2414: begin digit0<=FOUR; digit1<=ONE; digit2<=FOUR; digit3<=TWO; end
      16'd2415: begin digit0<=FIVE; digit1<=ONE; digit2<=FOUR; digit3<=TWO; end
      16'd2416: begin digit0<=SIX; digit1<=ONE; digit2<=FOUR; digit3<=TWO; end
      16'd2417: begin digit0<=SEVEN; digit1<=ONE; digit2<=FOUR; digit3<=TWO; end
      16'd2418: begin digit0<=EIGHT; digit1<=ONE; digit2<=FOUR; digit3<=TWO; end
      16'd2419: begin digit0<=NINE; digit1<=ONE; digit2<=FOUR; digit3<=TWO; end
      16'd2420: begin digit0<=ZERO; digit1<=TWO; digit2<=FOUR; digit3<=TWO; end
      16'd2421: begin digit0<=ONE; digit1<=TWO; digit2<=FOUR; digit3<=TWO; end
      16'd2422: begin digit0<=TWO; digit1<=TWO; digit2<=FOUR; digit3<=TWO; end
      16'd2423: begin digit0<=THREE; digit1<=TWO; digit2<=FOUR; digit3<=TWO; end
      16'd2424: begin digit0<=FOUR; digit1<=TWO; digit2<=FOUR; digit3<=TWO; end
      16'd2425: begin digit0<=FIVE; digit1<=TWO; digit2<=FOUR; digit3<=TWO; end
      16'd2426: begin digit0<=SIX; digit1<=TWO; digit2<=FOUR; digit3<=TWO; end
      16'd2427: begin digit0<=SEVEN; digit1<=TWO; digit2<=FOUR; digit3<=TWO; end
      16'd2428: begin digit0<=EIGHT; digit1<=TWO; digit2<=FOUR; digit3<=TWO; end
      16'd2429: begin digit0<=NINE; digit1<=TWO; digit2<=FOUR; digit3<=TWO; end
      16'd2430: begin digit0<=ZERO; digit1<=THREE; digit2<=FOUR; digit3<=TWO; end
      16'd2431: begin digit0<=ONE; digit1<=THREE; digit2<=FOUR; digit3<=TWO; end
      16'd2432: begin digit0<=TWO; digit1<=THREE; digit2<=FOUR; digit3<=TWO; end
      16'd2433: begin digit0<=THREE; digit1<=THREE; digit2<=FOUR; digit3<=TWO; end
      16'd2434: begin digit0<=FOUR; digit1<=THREE; digit2<=FOUR; digit3<=TWO; end
      16'd2435: begin digit0<=FIVE; digit1<=THREE; digit2<=FOUR; digit3<=TWO; end
      16'd2436: begin digit0<=SIX; digit1<=THREE; digit2<=FOUR; digit3<=TWO; end
      16'd2437: begin digit0<=SEVEN; digit1<=THREE; digit2<=FOUR; digit3<=TWO; end
      16'd2438: begin digit0<=EIGHT; digit1<=THREE; digit2<=FOUR; digit3<=TWO; end
      16'd2439: begin digit0<=NINE; digit1<=THREE; digit2<=FOUR; digit3<=TWO; end
      16'd2440: begin digit0<=ZERO; digit1<=FOUR; digit2<=FOUR; digit3<=TWO; end
      16'd2441: begin digit0<=ONE; digit1<=FOUR; digit2<=FOUR; digit3<=TWO; end
      16'd2442: begin digit0<=TWO; digit1<=FOUR; digit2<=FOUR; digit3<=TWO; end
      16'd2443: begin digit0<=THREE; digit1<=FOUR; digit2<=FOUR; digit3<=TWO; end
      16'd2444: begin digit0<=FOUR; digit1<=FOUR; digit2<=FOUR; digit3<=TWO; end
      16'd2445: begin digit0<=FIVE; digit1<=FOUR; digit2<=FOUR; digit3<=TWO; end
      16'd2446: begin digit0<=SIX; digit1<=FOUR; digit2<=FOUR; digit3<=TWO; end
      16'd2447: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FOUR; digit3<=TWO; end
      16'd2448: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FOUR; digit3<=TWO; end
      16'd2449: begin digit0<=NINE; digit1<=FOUR; digit2<=FOUR; digit3<=TWO; end
      16'd2450: begin digit0<=ZERO; digit1<=FIVE; digit2<=FOUR; digit3<=TWO; end
      16'd2451: begin digit0<=ONE; digit1<=FIVE; digit2<=FOUR; digit3<=TWO; end
      16'd2452: begin digit0<=TWO; digit1<=FIVE; digit2<=FOUR; digit3<=TWO; end
      16'd2453: begin digit0<=THREE; digit1<=FIVE; digit2<=FOUR; digit3<=TWO; end
      16'd2454: begin digit0<=FOUR; digit1<=FIVE; digit2<=FOUR; digit3<=TWO; end
      16'd2455: begin digit0<=FIVE; digit1<=FIVE; digit2<=FOUR; digit3<=TWO; end
      16'd2456: begin digit0<=SIX; digit1<=FIVE; digit2<=FOUR; digit3<=TWO; end
      16'd2457: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FOUR; digit3<=TWO; end
      16'd2458: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FOUR; digit3<=TWO; end
      16'd2459: begin digit0<=NINE; digit1<=FIVE; digit2<=FOUR; digit3<=TWO; end
      16'd2460: begin digit0<=ZERO; digit1<=SIX; digit2<=FOUR; digit3<=TWO; end
      16'd2461: begin digit0<=ONE; digit1<=SIX; digit2<=FOUR; digit3<=TWO; end
      16'd2462: begin digit0<=TWO; digit1<=SIX; digit2<=FOUR; digit3<=TWO; end
      16'd2463: begin digit0<=THREE; digit1<=SIX; digit2<=FOUR; digit3<=TWO; end
      16'd2464: begin digit0<=FOUR; digit1<=SIX; digit2<=FOUR; digit3<=TWO; end
      16'd2465: begin digit0<=FIVE; digit1<=SIX; digit2<=FOUR; digit3<=TWO; end
      16'd2466: begin digit0<=SIX; digit1<=SIX; digit2<=FOUR; digit3<=TWO; end
      16'd2467: begin digit0<=SEVEN; digit1<=SIX; digit2<=FOUR; digit3<=TWO; end
      16'd2468: begin digit0<=EIGHT; digit1<=SIX; digit2<=FOUR; digit3<=TWO; end
      16'd2469: begin digit0<=NINE; digit1<=SIX; digit2<=FOUR; digit3<=TWO; end
      16'd2470: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FOUR; digit3<=TWO; end
      16'd2471: begin digit0<=ONE; digit1<=SEVEN; digit2<=FOUR; digit3<=TWO; end
      16'd2472: begin digit0<=TWO; digit1<=SEVEN; digit2<=FOUR; digit3<=TWO; end
      16'd2473: begin digit0<=THREE; digit1<=SEVEN; digit2<=FOUR; digit3<=TWO; end
      16'd2474: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FOUR; digit3<=TWO; end
      16'd2475: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FOUR; digit3<=TWO; end
      16'd2476: begin digit0<=SIX; digit1<=SEVEN; digit2<=FOUR; digit3<=TWO; end
      16'd2477: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FOUR; digit3<=TWO; end
      16'd2478: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FOUR; digit3<=TWO; end
      16'd2479: begin digit0<=NINE; digit1<=SEVEN; digit2<=FOUR; digit3<=TWO; end
      16'd2480: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=TWO; end
      16'd2481: begin digit0<=ONE; digit1<=EIGHT; digit2<=FOUR; digit3<=TWO; end
      16'd2482: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=TWO; end
      16'd2483: begin digit0<=THREE; digit1<=EIGHT; digit2<=FOUR; digit3<=TWO; end
      16'd2484: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FOUR; digit3<=TWO; end
      16'd2485: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FOUR; digit3<=TWO; end
      16'd2486: begin digit0<=SIX; digit1<=EIGHT; digit2<=FOUR; digit3<=TWO; end
      16'd2487: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FOUR; digit3<=TWO; end
      16'd2488: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FOUR; digit3<=TWO; end
      16'd2489: begin digit0<=NINE; digit1<=EIGHT; digit2<=FOUR; digit3<=TWO; end
      16'd2490: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=TWO; end
      16'd2491: begin digit0<=ONE; digit1<=NINE; digit2<=FOUR; digit3<=TWO; end
      16'd2492: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=TWO; end
      16'd2493: begin digit0<=THREE; digit1<=NINE; digit2<=FOUR; digit3<=TWO; end
      16'd2494: begin digit0<=FOUR; digit1<=NINE; digit2<=FOUR; digit3<=TWO; end
      16'd2495: begin digit0<=FIVE; digit1<=NINE; digit2<=FOUR; digit3<=TWO; end
      16'd2496: begin digit0<=SIX; digit1<=NINE; digit2<=FOUR; digit3<=TWO; end
      16'd2497: begin digit0<=SEVEN; digit1<=NINE; digit2<=FOUR; digit3<=TWO; end
      16'd2498: begin digit0<=EIGHT; digit1<=NINE; digit2<=FOUR; digit3<=TWO; end
      16'd2499: begin digit0<=NINE; digit1<=NINE; digit2<=FOUR; digit3<=TWO; end
	  16'd2500: begin digit0<=ZERO; digit1<=ZERO; digit2<=FIVE; digit3<=TWO; end
      16'd2501: begin digit0<=ONE; digit1<=ZERO; digit2<=FIVE; digit3<=TWO; end
      16'd2502: begin digit0<=TWO; digit1<=ZERO; digit2<=FIVE; digit3<=TWO; end
      16'd2503: begin digit0<=THREE; digit1<=ZERO; digit2<=FIVE; digit3<=TWO; end
      16'd2504: begin digit0<=FOUR; digit1<=ZERO; digit2<=FIVE; digit3<=TWO; end
      16'd2505: begin digit0<=FIVE; digit1<=ZERO; digit2<=FIVE; digit3<=TWO; end
      16'd2506: begin digit0<=SIX; digit1<=ZERO; digit2<=FIVE; digit3<=TWO; end
      16'd2507: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FIVE; digit3<=TWO; end
      16'd2508: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FIVE; digit3<=TWO; end
      16'd2509: begin digit0<=NINE; digit1<=ZERO; digit2<=FIVE; digit3<=TWO; end
      16'd2510: begin digit0<=ZERO; digit1<=ONE; digit2<=FIVE; digit3<=TWO; end
      16'd2511: begin digit0<=ONE; digit1<=ONE; digit2<=FIVE; digit3<=TWO; end
      16'd2512: begin digit0<=TWO; digit1<=ONE; digit2<=FIVE; digit3<=TWO; end
      16'd2513: begin digit0<=THREE; digit1<=ONE; digit2<=FIVE; digit3<=TWO; end
      16'd2514: begin digit0<=FOUR; digit1<=ONE; digit2<=FIVE; digit3<=TWO; end
      16'd2515: begin digit0<=FIVE; digit1<=ONE; digit2<=FIVE; digit3<=TWO; end
      16'd2516: begin digit0<=SIX; digit1<=ONE; digit2<=FIVE; digit3<=TWO; end
      16'd2517: begin digit0<=SEVEN; digit1<=ONE; digit2<=FIVE; digit3<=TWO; end
      16'd2518: begin digit0<=EIGHT; digit1<=ONE; digit2<=FIVE; digit3<=TWO; end
      16'd2519: begin digit0<=NINE; digit1<=ONE; digit2<=FIVE; digit3<=TWO; end
      16'd2520: begin digit0<=ZERO; digit1<=TWO; digit2<=FIVE; digit3<=TWO; end
      16'd2521: begin digit0<=ONE; digit1<=TWO; digit2<=FIVE; digit3<=TWO; end
      16'd2522: begin digit0<=TWO; digit1<=TWO; digit2<=FIVE; digit3<=TWO; end
      16'd2523: begin digit0<=THREE; digit1<=TWO; digit2<=FIVE; digit3<=TWO; end
      16'd2524: begin digit0<=FOUR; digit1<=TWO; digit2<=FIVE; digit3<=TWO; end
      16'd2525: begin digit0<=FIVE; digit1<=TWO; digit2<=FIVE; digit3<=TWO; end
      16'd2526: begin digit0<=SIX; digit1<=TWO; digit2<=FIVE; digit3<=TWO; end
      16'd2527: begin digit0<=SEVEN; digit1<=TWO; digit2<=FIVE; digit3<=TWO; end
      16'd2528: begin digit0<=EIGHT; digit1<=TWO; digit2<=FIVE; digit3<=TWO; end
      16'd2529: begin digit0<=NINE; digit1<=TWO; digit2<=FIVE; digit3<=TWO; end
      16'd2530: begin digit0<=ZERO; digit1<=THREE; digit2<=FIVE; digit3<=TWO; end
      16'd2531: begin digit0<=ONE; digit1<=THREE; digit2<=FIVE; digit3<=TWO; end
      16'd2532: begin digit0<=TWO; digit1<=THREE; digit2<=FIVE; digit3<=TWO; end
      16'd2533: begin digit0<=THREE; digit1<=THREE; digit2<=FIVE; digit3<=TWO; end
      16'd2534: begin digit0<=FOUR; digit1<=THREE; digit2<=FIVE; digit3<=TWO; end
      16'd2535: begin digit0<=FIVE; digit1<=THREE; digit2<=FIVE; digit3<=TWO; end
      16'd2536: begin digit0<=SIX; digit1<=THREE; digit2<=FIVE; digit3<=TWO; end
      16'd2537: begin digit0<=SEVEN; digit1<=THREE; digit2<=FIVE; digit3<=TWO; end
      16'd2538: begin digit0<=EIGHT; digit1<=THREE; digit2<=FIVE; digit3<=TWO; end
      16'd2539: begin digit0<=NINE; digit1<=THREE; digit2<=FIVE; digit3<=TWO; end
      16'd2540: begin digit0<=ZERO; digit1<=FOUR; digit2<=FIVE; digit3<=TWO; end
      16'd2541: begin digit0<=ONE; digit1<=FOUR; digit2<=FIVE; digit3<=TWO; end
      16'd2542: begin digit0<=TWO; digit1<=FOUR; digit2<=FIVE; digit3<=TWO; end
      16'd2543: begin digit0<=THREE; digit1<=FOUR; digit2<=FIVE; digit3<=TWO; end
      16'd2544: begin digit0<=FOUR; digit1<=FOUR; digit2<=FIVE; digit3<=TWO; end
      16'd2545: begin digit0<=FIVE; digit1<=FOUR; digit2<=FIVE; digit3<=TWO; end
      16'd2546: begin digit0<=SIX; digit1<=FOUR; digit2<=FIVE; digit3<=TWO; end
      16'd2547: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FIVE; digit3<=TWO; end
      16'd2548: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FIVE; digit3<=TWO; end
      16'd2549: begin digit0<=NINE; digit1<=FOUR; digit2<=FIVE; digit3<=TWO; end
      16'd2550: begin digit0<=ZERO; digit1<=FIVE; digit2<=FIVE; digit3<=TWO; end
      16'd2551: begin digit0<=ONE; digit1<=FIVE; digit2<=FIVE; digit3<=TWO; end
      16'd2552: begin digit0<=TWO; digit1<=FIVE; digit2<=FIVE; digit3<=TWO; end
      16'd2553: begin digit0<=THREE; digit1<=FIVE; digit2<=FIVE; digit3<=TWO; end
      16'd2554: begin digit0<=FOUR; digit1<=FIVE; digit2<=FIVE; digit3<=TWO; end
      16'd2555: begin digit0<=FIVE; digit1<=FIVE; digit2<=FIVE; digit3<=TWO; end
      16'd2556: begin digit0<=SIX; digit1<=FIVE; digit2<=FIVE; digit3<=TWO; end
      16'd2557: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FIVE; digit3<=TWO; end
      16'd2558: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FIVE; digit3<=TWO; end
      16'd2559: begin digit0<=NINE; digit1<=FIVE; digit2<=FIVE; digit3<=TWO; end
      16'd2560: begin digit0<=ZERO; digit1<=SIX; digit2<=FIVE; digit3<=TWO; end
      16'd2561: begin digit0<=ONE; digit1<=SIX; digit2<=FIVE; digit3<=TWO; end
      16'd2562: begin digit0<=TWO; digit1<=SIX; digit2<=FIVE; digit3<=TWO; end
      16'd2563: begin digit0<=THREE; digit1<=SIX; digit2<=FIVE; digit3<=TWO; end
      16'd2564: begin digit0<=FOUR; digit1<=SIX; digit2<=FIVE; digit3<=TWO; end
      16'd2565: begin digit0<=FIVE; digit1<=SIX; digit2<=FIVE; digit3<=TWO; end
      16'd2566: begin digit0<=SIX; digit1<=SIX; digit2<=FIVE; digit3<=TWO; end
      16'd2567: begin digit0<=SEVEN; digit1<=SIX; digit2<=FIVE; digit3<=TWO; end
      16'd2568: begin digit0<=EIGHT; digit1<=SIX; digit2<=FIVE; digit3<=TWO; end
      16'd2569: begin digit0<=NINE; digit1<=SIX; digit2<=FIVE; digit3<=TWO; end
      16'd2570: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FIVE; digit3<=TWO; end
      16'd2571: begin digit0<=ONE; digit1<=SEVEN; digit2<=FIVE; digit3<=TWO; end
      16'd2572: begin digit0<=TWO; digit1<=SEVEN; digit2<=FIVE; digit3<=TWO; end
      16'd2573: begin digit0<=THREE; digit1<=SEVEN; digit2<=FIVE; digit3<=TWO; end
      16'd2574: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FIVE; digit3<=TWO; end
      16'd2575: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FIVE; digit3<=TWO; end
      16'd2576: begin digit0<=SIX; digit1<=SEVEN; digit2<=FIVE; digit3<=TWO; end
      16'd2577: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FIVE; digit3<=TWO; end
      16'd2578: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FIVE; digit3<=TWO; end
      16'd2579: begin digit0<=NINE; digit1<=SEVEN; digit2<=FIVE; digit3<=TWO; end
      16'd2580: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=TWO; end
      16'd2581: begin digit0<=ONE; digit1<=EIGHT; digit2<=FIVE; digit3<=TWO; end
      16'd2582: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=TWO; end
      16'd2583: begin digit0<=THREE; digit1<=EIGHT; digit2<=FIVE; digit3<=TWO; end
      16'd2584: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FIVE; digit3<=TWO; end
      16'd2585: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FIVE; digit3<=TWO; end
      16'd2586: begin digit0<=SIX; digit1<=EIGHT; digit2<=FIVE; digit3<=TWO; end
      16'd2587: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FIVE; digit3<=TWO; end
      16'd2588: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FIVE; digit3<=TWO; end
      16'd2589: begin digit0<=NINE; digit1<=EIGHT; digit2<=FIVE; digit3<=TWO; end
      16'd2590: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=TWO; end
      16'd2591: begin digit0<=ONE; digit1<=NINE; digit2<=FIVE; digit3<=TWO; end
      16'd2592: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=TWO; end
      16'd2593: begin digit0<=THREE; digit1<=NINE; digit2<=FIVE; digit3<=TWO; end
      16'd2594: begin digit0<=FOUR; digit1<=NINE; digit2<=FIVE; digit3<=TWO; end
      16'd2595: begin digit0<=FIVE; digit1<=NINE; digit2<=FIVE; digit3<=TWO; end
      16'd2596: begin digit0<=SIX; digit1<=NINE; digit2<=FIVE; digit3<=TWO; end
      16'd2597: begin digit0<=SEVEN; digit1<=NINE; digit2<=FIVE; digit3<=TWO; end
      16'd2598: begin digit0<=EIGHT; digit1<=NINE; digit2<=FIVE; digit3<=TWO; end
      16'd2599: begin digit0<=NINE; digit1<=NINE; digit2<=FIVE; digit3<=TWO; end
	  16'd2600: begin digit0<=ZERO; digit1<=ZERO; digit2<=SIX; digit3<=TWO; end
      16'd2601: begin digit0<=ONE; digit1<=ZERO; digit2<=SIX; digit3<=TWO; end
      16'd2602: begin digit0<=TWO; digit1<=ZERO; digit2<=SIX; digit3<=TWO; end
      16'd2603: begin digit0<=THREE; digit1<=ZERO; digit2<=SIX; digit3<=TWO; end
      16'd2604: begin digit0<=FOUR; digit1<=ZERO; digit2<=SIX; digit3<=TWO; end
      16'd2605: begin digit0<=FIVE; digit1<=ZERO; digit2<=SIX; digit3<=TWO; end
      16'd2606: begin digit0<=SIX; digit1<=ZERO; digit2<=SIX; digit3<=TWO; end
      16'd2607: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SIX; digit3<=TWO; end
      16'd2608: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SIX; digit3<=TWO; end
      16'd2609: begin digit0<=NINE; digit1<=ZERO; digit2<=SIX; digit3<=TWO; end
      16'd2610: begin digit0<=ZERO; digit1<=ONE; digit2<=SIX; digit3<=TWO; end
      16'd2611: begin digit0<=ONE; digit1<=ONE; digit2<=SIX; digit3<=TWO; end
      16'd2612: begin digit0<=TWO; digit1<=ONE; digit2<=SIX; digit3<=TWO; end
      16'd2613: begin digit0<=THREE; digit1<=ONE; digit2<=SIX; digit3<=TWO; end
      16'd2614: begin digit0<=FOUR; digit1<=ONE; digit2<=SIX; digit3<=TWO; end
      16'd2615: begin digit0<=FIVE; digit1<=ONE; digit2<=SIX; digit3<=TWO; end
      16'd2616: begin digit0<=SIX; digit1<=ONE; digit2<=SIX; digit3<=TWO; end
      16'd2617: begin digit0<=SEVEN; digit1<=ONE; digit2<=SIX; digit3<=TWO; end
      16'd2618: begin digit0<=EIGHT; digit1<=ONE; digit2<=SIX; digit3<=TWO; end
      16'd2619: begin digit0<=NINE; digit1<=ONE; digit2<=SIX; digit3<=TWO; end
      16'd2620: begin digit0<=ZERO; digit1<=TWO; digit2<=SIX; digit3<=TWO; end
      16'd2621: begin digit0<=ONE; digit1<=TWO; digit2<=SIX; digit3<=TWO; end
      16'd2622: begin digit0<=TWO; digit1<=TWO; digit2<=SIX; digit3<=TWO; end
      16'd2623: begin digit0<=THREE; digit1<=TWO; digit2<=SIX; digit3<=TWO; end
      16'd2624: begin digit0<=FOUR; digit1<=TWO; digit2<=SIX; digit3<=TWO; end
      16'd2625: begin digit0<=FIVE; digit1<=TWO; digit2<=SIX; digit3<=TWO; end
      16'd2626: begin digit0<=SIX; digit1<=TWO; digit2<=SIX; digit3<=TWO; end
      16'd2627: begin digit0<=SEVEN; digit1<=TWO; digit2<=SIX; digit3<=TWO; end
      16'd2628: begin digit0<=EIGHT; digit1<=TWO; digit2<=SIX; digit3<=TWO; end
      16'd2629: begin digit0<=NINE; digit1<=TWO; digit2<=SIX; digit3<=TWO; end
      16'd2630: begin digit0<=ZERO; digit1<=THREE; digit2<=SIX; digit3<=TWO; end
      16'd2631: begin digit0<=ONE; digit1<=THREE; digit2<=SIX; digit3<=TWO; end
      16'd2632: begin digit0<=TWO; digit1<=THREE; digit2<=SIX; digit3<=TWO; end
      16'd2633: begin digit0<=THREE; digit1<=THREE; digit2<=SIX; digit3<=TWO; end
      16'd2634: begin digit0<=FOUR; digit1<=THREE; digit2<=SIX; digit3<=TWO; end
      16'd2635: begin digit0<=FIVE; digit1<=THREE; digit2<=SIX; digit3<=TWO; end
      16'd2636: begin digit0<=SIX; digit1<=THREE; digit2<=SIX; digit3<=TWO; end
      16'd2637: begin digit0<=SEVEN; digit1<=THREE; digit2<=SIX; digit3<=TWO; end
      16'd2638: begin digit0<=EIGHT; digit1<=THREE; digit2<=SIX; digit3<=TWO; end
      16'd2639: begin digit0<=NINE; digit1<=THREE; digit2<=SIX; digit3<=TWO; end
      16'd2640: begin digit0<=ZERO; digit1<=FOUR; digit2<=SIX; digit3<=TWO; end
      16'd2641: begin digit0<=ONE; digit1<=FOUR; digit2<=SIX; digit3<=TWO; end
      16'd2642: begin digit0<=TWO; digit1<=FOUR; digit2<=SIX; digit3<=TWO; end
      16'd2643: begin digit0<=THREE; digit1<=FOUR; digit2<=SIX; digit3<=TWO; end
      16'd2644: begin digit0<=FOUR; digit1<=FOUR; digit2<=SIX; digit3<=TWO; end
      16'd2645: begin digit0<=FIVE; digit1<=FOUR; digit2<=SIX; digit3<=TWO; end
      16'd2646: begin digit0<=SIX; digit1<=FOUR; digit2<=SIX; digit3<=TWO; end
      16'd2647: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SIX; digit3<=TWO; end
      16'd2648: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SIX; digit3<=TWO; end
      16'd2649: begin digit0<=NINE; digit1<=FOUR; digit2<=SIX; digit3<=TWO; end
      16'd2650: begin digit0<=ZERO; digit1<=FIVE; digit2<=SIX; digit3<=TWO; end
      16'd2651: begin digit0<=ONE; digit1<=FIVE; digit2<=SIX; digit3<=TWO; end
      16'd2652: begin digit0<=TWO; digit1<=FIVE; digit2<=SIX; digit3<=TWO; end
      16'd2653: begin digit0<=THREE; digit1<=FIVE; digit2<=SIX; digit3<=TWO; end
      16'd2654: begin digit0<=FOUR; digit1<=FIVE; digit2<=SIX; digit3<=TWO; end
      16'd2655: begin digit0<=FIVE; digit1<=FIVE; digit2<=SIX; digit3<=TWO; end
      16'd2656: begin digit0<=SIX; digit1<=FIVE; digit2<=SIX; digit3<=TWO; end
      16'd2657: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SIX; digit3<=TWO; end
      16'd2658: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SIX; digit3<=TWO; end
      16'd2659: begin digit0<=NINE; digit1<=FIVE; digit2<=SIX; digit3<=TWO; end
      16'd2660: begin digit0<=ZERO; digit1<=SIX; digit2<=SIX; digit3<=TWO; end
      16'd2661: begin digit0<=ONE; digit1<=SIX; digit2<=SIX; digit3<=TWO; end
      16'd2662: begin digit0<=TWO; digit1<=SIX; digit2<=SIX; digit3<=TWO; end
      16'd2663: begin digit0<=THREE; digit1<=SIX; digit2<=SIX; digit3<=TWO; end
      16'd2664: begin digit0<=FOUR; digit1<=SIX; digit2<=SIX; digit3<=TWO; end
      16'd2665: begin digit0<=FIVE; digit1<=SIX; digit2<=SIX; digit3<=TWO; end
      16'd2666: begin digit0<=SIX; digit1<=SIX; digit2<=SIX; digit3<=TWO; end
      16'd2667: begin digit0<=SEVEN; digit1<=SIX; digit2<=SIX; digit3<=TWO; end
      16'd2668: begin digit0<=EIGHT; digit1<=SIX; digit2<=SIX; digit3<=TWO; end
      16'd2669: begin digit0<=NINE; digit1<=SIX; digit2<=SIX; digit3<=TWO; end
      16'd2670: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SIX; digit3<=TWO; end
      16'd2671: begin digit0<=ONE; digit1<=SEVEN; digit2<=SIX; digit3<=TWO; end
      16'd2672: begin digit0<=TWO; digit1<=SEVEN; digit2<=SIX; digit3<=TWO; end
      16'd2673: begin digit0<=THREE; digit1<=SEVEN; digit2<=SIX; digit3<=TWO; end
      16'd2674: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SIX; digit3<=TWO; end
      16'd2675: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SIX; digit3<=TWO; end
      16'd2676: begin digit0<=SIX; digit1<=SEVEN; digit2<=SIX; digit3<=TWO; end
      16'd2677: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SIX; digit3<=TWO; end
      16'd2678: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SIX; digit3<=TWO; end
      16'd2679: begin digit0<=NINE; digit1<=SEVEN; digit2<=SIX; digit3<=TWO; end
      16'd2680: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=TWO; end
      16'd2681: begin digit0<=ONE; digit1<=EIGHT; digit2<=SIX; digit3<=TWO; end
      16'd2682: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=TWO; end
      16'd2683: begin digit0<=THREE; digit1<=EIGHT; digit2<=SIX; digit3<=TWO; end
      16'd2684: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SIX; digit3<=TWO; end
      16'd2685: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SIX; digit3<=TWO; end
      16'd2686: begin digit0<=SIX; digit1<=EIGHT; digit2<=SIX; digit3<=TWO; end
      16'd2687: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SIX; digit3<=TWO; end
      16'd2688: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SIX; digit3<=TWO; end
      16'd2689: begin digit0<=NINE; digit1<=EIGHT; digit2<=SIX; digit3<=TWO; end
      16'd2690: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=TWO; end
      16'd2691: begin digit0<=ONE; digit1<=NINE; digit2<=SIX; digit3<=TWO; end
      16'd2692: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=TWO; end
      16'd2693: begin digit0<=THREE; digit1<=NINE; digit2<=SIX; digit3<=TWO; end
      16'd2694: begin digit0<=FOUR; digit1<=NINE; digit2<=SIX; digit3<=TWO; end
      16'd2695: begin digit0<=FIVE; digit1<=NINE; digit2<=SIX; digit3<=TWO; end
      16'd2696: begin digit0<=SIX; digit1<=NINE; digit2<=SIX; digit3<=TWO; end
      16'd2697: begin digit0<=SEVEN; digit1<=NINE; digit2<=SIX; digit3<=TWO; end
      16'd2698: begin digit0<=EIGHT; digit1<=NINE; digit2<=SIX; digit3<=TWO; end
      16'd2699: begin digit0<=NINE; digit1<=NINE; digit2<=SIX; digit3<=TWO; end
	  16'd2700: begin digit0<=ZERO; digit1<=ZERO; digit2<=SEVEN; digit3<=TWO; end
      16'd2701: begin digit0<=ONE; digit1<=ZERO; digit2<=SEVEN; digit3<=TWO; end
      16'd2702: begin digit0<=TWO; digit1<=ZERO; digit2<=SEVEN; digit3<=TWO; end
      16'd2703: begin digit0<=THREE; digit1<=ZERO; digit2<=SEVEN; digit3<=TWO; end
      16'd2704: begin digit0<=FOUR; digit1<=ZERO; digit2<=SEVEN; digit3<=TWO; end
      16'd2705: begin digit0<=FIVE; digit1<=ZERO; digit2<=SEVEN; digit3<=TWO; end
      16'd2706: begin digit0<=SIX; digit1<=ZERO; digit2<=SEVEN; digit3<=TWO; end
      16'd2707: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SEVEN; digit3<=TWO; end
      16'd2708: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SEVEN; digit3<=TWO; end
      16'd2709: begin digit0<=NINE; digit1<=ZERO; digit2<=SEVEN; digit3<=TWO; end
      16'd2710: begin digit0<=ZERO; digit1<=ONE; digit2<=SEVEN; digit3<=TWO; end
      16'd2711: begin digit0<=ONE; digit1<=ONE; digit2<=SEVEN; digit3<=TWO; end
      16'd2712: begin digit0<=TWO; digit1<=ONE; digit2<=SEVEN; digit3<=TWO; end
      16'd2713: begin digit0<=THREE; digit1<=ONE; digit2<=SEVEN; digit3<=TWO; end
      16'd2714: begin digit0<=FOUR; digit1<=ONE; digit2<=SEVEN; digit3<=TWO; end
      16'd2715: begin digit0<=FIVE; digit1<=ONE; digit2<=SEVEN; digit3<=TWO; end
      16'd2716: begin digit0<=SIX; digit1<=ONE; digit2<=SEVEN; digit3<=TWO; end
      16'd2717: begin digit0<=SEVEN; digit1<=ONE; digit2<=SEVEN; digit3<=TWO; end
      16'd2718: begin digit0<=EIGHT; digit1<=ONE; digit2<=SEVEN; digit3<=TWO; end
      16'd2719: begin digit0<=NINE; digit1<=ONE; digit2<=SEVEN; digit3<=TWO; end
      16'd2720: begin digit0<=ZERO; digit1<=TWO; digit2<=SEVEN; digit3<=TWO; end
      16'd2721: begin digit0<=ONE; digit1<=TWO; digit2<=SEVEN; digit3<=TWO; end
      16'd2722: begin digit0<=TWO; digit1<=TWO; digit2<=SEVEN; digit3<=TWO; end
      16'd2723: begin digit0<=THREE; digit1<=TWO; digit2<=SEVEN; digit3<=TWO; end
      16'd2724: begin digit0<=FOUR; digit1<=TWO; digit2<=SEVEN; digit3<=TWO; end
      16'd2725: begin digit0<=FIVE; digit1<=TWO; digit2<=SEVEN; digit3<=TWO; end
      16'd2726: begin digit0<=SIX; digit1<=TWO; digit2<=SEVEN; digit3<=TWO; end
      16'd2727: begin digit0<=SEVEN; digit1<=TWO; digit2<=SEVEN; digit3<=TWO; end
      16'd2728: begin digit0<=EIGHT; digit1<=TWO; digit2<=SEVEN; digit3<=TWO; end
      16'd2729: begin digit0<=NINE; digit1<=TWO; digit2<=SEVEN; digit3<=TWO; end
      16'd2730: begin digit0<=ZERO; digit1<=THREE; digit2<=SEVEN; digit3<=TWO; end
      16'd2731: begin digit0<=ONE; digit1<=THREE; digit2<=SEVEN; digit3<=TWO; end
      16'd2732: begin digit0<=TWO; digit1<=THREE; digit2<=SEVEN; digit3<=TWO; end
      16'd2733: begin digit0<=THREE; digit1<=THREE; digit2<=SEVEN; digit3<=TWO; end
      16'd2734: begin digit0<=FOUR; digit1<=THREE; digit2<=SEVEN; digit3<=TWO; end
      16'd2735: begin digit0<=FIVE; digit1<=THREE; digit2<=SEVEN; digit3<=TWO; end
      16'd2736: begin digit0<=SIX; digit1<=THREE; digit2<=SEVEN; digit3<=TWO; end
      16'd2737: begin digit0<=SEVEN; digit1<=THREE; digit2<=SEVEN; digit3<=TWO; end
      16'd2738: begin digit0<=EIGHT; digit1<=THREE; digit2<=SEVEN; digit3<=TWO; end
      16'd2739: begin digit0<=NINE; digit1<=THREE; digit2<=SEVEN; digit3<=TWO; end
      16'd2740: begin digit0<=ZERO; digit1<=FOUR; digit2<=SEVEN; digit3<=TWO; end
      16'd2741: begin digit0<=ONE; digit1<=FOUR; digit2<=SEVEN; digit3<=TWO; end
      16'd2742: begin digit0<=TWO; digit1<=FOUR; digit2<=SEVEN; digit3<=TWO; end
      16'd2743: begin digit0<=THREE; digit1<=FOUR; digit2<=SEVEN; digit3<=TWO; end
      16'd2744: begin digit0<=FOUR; digit1<=FOUR; digit2<=SEVEN; digit3<=TWO; end
      16'd2745: begin digit0<=FIVE; digit1<=FOUR; digit2<=SEVEN; digit3<=TWO; end
      16'd2746: begin digit0<=SIX; digit1<=FOUR; digit2<=SEVEN; digit3<=TWO; end
      16'd2747: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SEVEN; digit3<=TWO; end
      16'd2748: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SEVEN; digit3<=TWO; end
      16'd2749: begin digit0<=NINE; digit1<=FOUR; digit2<=SEVEN; digit3<=TWO; end
      16'd2750: begin digit0<=ZERO; digit1<=FIVE; digit2<=SEVEN; digit3<=TWO; end
      16'd2751: begin digit0<=ONE; digit1<=FIVE; digit2<=SEVEN; digit3<=TWO; end
      16'd2752: begin digit0<=TWO; digit1<=FIVE; digit2<=SEVEN; digit3<=TWO; end
      16'd2753: begin digit0<=THREE; digit1<=FIVE; digit2<=SEVEN; digit3<=TWO; end
      16'd2754: begin digit0<=FOUR; digit1<=FIVE; digit2<=SEVEN; digit3<=TWO; end
      16'd2755: begin digit0<=FIVE; digit1<=FIVE; digit2<=SEVEN; digit3<=TWO; end
      16'd2756: begin digit0<=SIX; digit1<=FIVE; digit2<=SEVEN; digit3<=TWO; end
      16'd2757: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SEVEN; digit3<=TWO; end
      16'd2758: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SEVEN; digit3<=TWO; end
      16'd2759: begin digit0<=NINE; digit1<=FIVE; digit2<=SEVEN; digit3<=TWO; end
      16'd2760: begin digit0<=ZERO; digit1<=SIX; digit2<=SEVEN; digit3<=TWO; end
      16'd2761: begin digit0<=ONE; digit1<=SIX; digit2<=SEVEN; digit3<=TWO; end
      16'd2762: begin digit0<=TWO; digit1<=SIX; digit2<=SEVEN; digit3<=TWO; end
      16'd2763: begin digit0<=THREE; digit1<=SIX; digit2<=SEVEN; digit3<=TWO; end
      16'd2764: begin digit0<=FOUR; digit1<=SIX; digit2<=SEVEN; digit3<=TWO; end
      16'd2765: begin digit0<=FIVE; digit1<=SIX; digit2<=SEVEN; digit3<=TWO; end
      16'd2766: begin digit0<=SIX; digit1<=SIX; digit2<=SEVEN; digit3<=TWO; end
      16'd2767: begin digit0<=SEVEN; digit1<=SIX; digit2<=SEVEN; digit3<=TWO; end
      16'd2768: begin digit0<=EIGHT; digit1<=SIX; digit2<=SEVEN; digit3<=TWO; end
      16'd2769: begin digit0<=NINE; digit1<=SIX; digit2<=SEVEN; digit3<=TWO; end
      16'd2770: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SEVEN; digit3<=TWO; end
      16'd2771: begin digit0<=ONE; digit1<=SEVEN; digit2<=SEVEN; digit3<=TWO; end
      16'd2772: begin digit0<=TWO; digit1<=SEVEN; digit2<=SEVEN; digit3<=TWO; end
      16'd2773: begin digit0<=THREE; digit1<=SEVEN; digit2<=SEVEN; digit3<=TWO; end
      16'd2774: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SEVEN; digit3<=TWO; end
      16'd2775: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SEVEN; digit3<=TWO; end
      16'd2776: begin digit0<=SIX; digit1<=SEVEN; digit2<=SEVEN; digit3<=TWO; end
      16'd2777: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SEVEN; digit3<=TWO; end
      16'd2778: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SEVEN; digit3<=TWO; end
      16'd2779: begin digit0<=NINE; digit1<=SEVEN; digit2<=SEVEN; digit3<=TWO; end
      16'd2780: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=TWO; end
      16'd2781: begin digit0<=ONE; digit1<=EIGHT; digit2<=SEVEN; digit3<=TWO; end
      16'd2782: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=TWO; end
      16'd2783: begin digit0<=THREE; digit1<=EIGHT; digit2<=SEVEN; digit3<=TWO; end
      16'd2784: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SEVEN; digit3<=TWO; end
      16'd2785: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SEVEN; digit3<=TWO; end
      16'd2786: begin digit0<=SIX; digit1<=EIGHT; digit2<=SEVEN; digit3<=TWO; end
      16'd2787: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SEVEN; digit3<=TWO; end
      16'd2788: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SEVEN; digit3<=TWO; end
      16'd2789: begin digit0<=NINE; digit1<=EIGHT; digit2<=SEVEN; digit3<=TWO; end
      16'd2790: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=TWO; end
      16'd2791: begin digit0<=ONE; digit1<=NINE; digit2<=SEVEN; digit3<=TWO; end
      16'd2792: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=TWO; end
      16'd2793: begin digit0<=THREE; digit1<=NINE; digit2<=SEVEN; digit3<=TWO; end
      16'd2794: begin digit0<=FOUR; digit1<=NINE; digit2<=SEVEN; digit3<=TWO; end
      16'd2795: begin digit0<=FIVE; digit1<=NINE; digit2<=SEVEN; digit3<=TWO; end
      16'd2796: begin digit0<=SIX; digit1<=NINE; digit2<=SEVEN; digit3<=TWO; end
      16'd2797: begin digit0<=SEVEN; digit1<=NINE; digit2<=SEVEN; digit3<=TWO; end
      16'd2798: begin digit0<=EIGHT; digit1<=NINE; digit2<=SEVEN; digit3<=TWO; end
      16'd2799: begin digit0<=NINE; digit1<=NINE; digit2<=SEVEN; digit3<=TWO; end
	  16'd2800: begin digit0<=ZERO; digit1<=ZERO; digit2<=EIGHT; digit3<=TWO; end
      16'd2801: begin digit0<=ONE; digit1<=ZERO; digit2<=EIGHT; digit3<=TWO; end
      16'd2802: begin digit0<=TWO; digit1<=ZERO; digit2<=EIGHT; digit3<=TWO; end
      16'd2803: begin digit0<=THREE; digit1<=ZERO; digit2<=EIGHT; digit3<=TWO; end
      16'd2804: begin digit0<=FOUR; digit1<=ZERO; digit2<=EIGHT; digit3<=TWO; end
      16'd2805: begin digit0<=FIVE; digit1<=ZERO; digit2<=EIGHT; digit3<=TWO; end
      16'd2806: begin digit0<=SIX; digit1<=ZERO; digit2<=EIGHT; digit3<=TWO; end
      16'd2807: begin digit0<=SEVEN; digit1<=ZERO; digit2<=EIGHT; digit3<=TWO; end
      16'd2808: begin digit0<=EIGHT; digit1<=ZERO; digit2<=EIGHT; digit3<=TWO; end
      16'd2809: begin digit0<=NINE; digit1<=ZERO; digit2<=EIGHT; digit3<=TWO; end
      16'd2810: begin digit0<=ZERO; digit1<=ONE; digit2<=EIGHT; digit3<=TWO; end
      16'd2811: begin digit0<=ONE; digit1<=ONE; digit2<=EIGHT; digit3<=TWO; end
      16'd2812: begin digit0<=TWO; digit1<=ONE; digit2<=EIGHT; digit3<=TWO; end
      16'd2813: begin digit0<=THREE; digit1<=ONE; digit2<=EIGHT; digit3<=TWO; end
      16'd2814: begin digit0<=FOUR; digit1<=ONE; digit2<=EIGHT; digit3<=TWO; end
      16'd2815: begin digit0<=FIVE; digit1<=ONE; digit2<=EIGHT; digit3<=TWO; end
      16'd2816: begin digit0<=SIX; digit1<=ONE; digit2<=EIGHT; digit3<=TWO; end
      16'd2817: begin digit0<=SEVEN; digit1<=ONE; digit2<=EIGHT; digit3<=TWO; end
      16'd2818: begin digit0<=EIGHT; digit1<=ONE; digit2<=EIGHT; digit3<=TWO; end
      16'd2819: begin digit0<=NINE; digit1<=ONE; digit2<=EIGHT; digit3<=TWO; end
      16'd2820: begin digit0<=ZERO; digit1<=TWO; digit2<=EIGHT; digit3<=TWO; end
      16'd2821: begin digit0<=ONE; digit1<=TWO; digit2<=EIGHT; digit3<=TWO; end
      16'd2822: begin digit0<=TWO; digit1<=TWO; digit2<=EIGHT; digit3<=TWO; end
      16'd2823: begin digit0<=THREE; digit1<=TWO; digit2<=EIGHT; digit3<=TWO; end
      16'd2824: begin digit0<=FOUR; digit1<=TWO; digit2<=EIGHT; digit3<=TWO; end
      16'd2825: begin digit0<=FIVE; digit1<=TWO; digit2<=EIGHT; digit3<=TWO; end
      16'd2826: begin digit0<=SIX; digit1<=TWO; digit2<=EIGHT; digit3<=TWO; end
      16'd2827: begin digit0<=SEVEN; digit1<=TWO; digit2<=EIGHT; digit3<=TWO; end
      16'd2828: begin digit0<=EIGHT; digit1<=TWO; digit2<=EIGHT; digit3<=TWO; end
      16'd2829: begin digit0<=NINE; digit1<=TWO; digit2<=EIGHT; digit3<=TWO; end
      16'd2830: begin digit0<=ZERO; digit1<=THREE; digit2<=EIGHT; digit3<=TWO; end
      16'd2831: begin digit0<=ONE; digit1<=THREE; digit2<=EIGHT; digit3<=TWO; end
      16'd2832: begin digit0<=TWO; digit1<=THREE; digit2<=EIGHT; digit3<=TWO; end
      16'd2833: begin digit0<=THREE; digit1<=THREE; digit2<=EIGHT; digit3<=TWO; end
      16'd2834: begin digit0<=FOUR; digit1<=THREE; digit2<=EIGHT; digit3<=TWO; end
      16'd2835: begin digit0<=FIVE; digit1<=THREE; digit2<=EIGHT; digit3<=TWO; end
      16'd2836: begin digit0<=SIX; digit1<=THREE; digit2<=EIGHT; digit3<=TWO; end
      16'd2837: begin digit0<=SEVEN; digit1<=THREE; digit2<=EIGHT; digit3<=TWO; end
      16'd2838: begin digit0<=EIGHT; digit1<=THREE; digit2<=EIGHT; digit3<=TWO; end
      16'd2839: begin digit0<=NINE; digit1<=THREE; digit2<=EIGHT; digit3<=TWO; end
      16'd2840: begin digit0<=ZERO; digit1<=FOUR; digit2<=EIGHT; digit3<=TWO; end
      16'd2841: begin digit0<=ONE; digit1<=FOUR; digit2<=EIGHT; digit3<=TWO; end
      16'd2842: begin digit0<=TWO; digit1<=FOUR; digit2<=EIGHT; digit3<=TWO; end
      16'd2843: begin digit0<=THREE; digit1<=FOUR; digit2<=EIGHT; digit3<=TWO; end
      16'd2844: begin digit0<=FOUR; digit1<=FOUR; digit2<=EIGHT; digit3<=TWO; end
      16'd2845: begin digit0<=FIVE; digit1<=FOUR; digit2<=EIGHT; digit3<=TWO; end
      16'd2846: begin digit0<=SIX; digit1<=FOUR; digit2<=EIGHT; digit3<=TWO; end
      16'd2847: begin digit0<=SEVEN; digit1<=FOUR; digit2<=EIGHT; digit3<=TWO; end
      16'd2848: begin digit0<=EIGHT; digit1<=FOUR; digit2<=EIGHT; digit3<=TWO; end
      16'd2849: begin digit0<=NINE; digit1<=FOUR; digit2<=EIGHT; digit3<=TWO; end
      16'd2850: begin digit0<=ZERO; digit1<=FIVE; digit2<=EIGHT; digit3<=TWO; end
      16'd2851: begin digit0<=ONE; digit1<=FIVE; digit2<=EIGHT; digit3<=TWO; end
      16'd2852: begin digit0<=TWO; digit1<=FIVE; digit2<=EIGHT; digit3<=TWO; end
      16'd2853: begin digit0<=THREE; digit1<=FIVE; digit2<=EIGHT; digit3<=TWO; end
      16'd2854: begin digit0<=FOUR; digit1<=FIVE; digit2<=EIGHT; digit3<=TWO; end
      16'd2855: begin digit0<=FIVE; digit1<=FIVE; digit2<=EIGHT; digit3<=TWO; end
      16'd2856: begin digit0<=SIX; digit1<=FIVE; digit2<=EIGHT; digit3<=TWO; end
      16'd2857: begin digit0<=SEVEN; digit1<=FIVE; digit2<=EIGHT; digit3<=TWO; end
      16'd2858: begin digit0<=EIGHT; digit1<=FIVE; digit2<=EIGHT; digit3<=TWO; end
      16'd2859: begin digit0<=NINE; digit1<=FIVE; digit2<=EIGHT; digit3<=TWO; end
      16'd2860: begin digit0<=ZERO; digit1<=SIX; digit2<=EIGHT; digit3<=TWO; end
      16'd2861: begin digit0<=ONE; digit1<=SIX; digit2<=EIGHT; digit3<=TWO; end
      16'd2862: begin digit0<=TWO; digit1<=SIX; digit2<=EIGHT; digit3<=TWO; end
      16'd2863: begin digit0<=THREE; digit1<=SIX; digit2<=EIGHT; digit3<=TWO; end
      16'd2864: begin digit0<=FOUR; digit1<=SIX; digit2<=EIGHT; digit3<=TWO; end
      16'd2865: begin digit0<=FIVE; digit1<=SIX; digit2<=EIGHT; digit3<=TWO; end
      16'd2866: begin digit0<=SIX; digit1<=SIX; digit2<=EIGHT; digit3<=TWO; end
      16'd2867: begin digit0<=SEVEN; digit1<=SIX; digit2<=EIGHT; digit3<=TWO; end
      16'd2868: begin digit0<=EIGHT; digit1<=SIX; digit2<=EIGHT; digit3<=TWO; end
      16'd2869: begin digit0<=NINE; digit1<=SIX; digit2<=EIGHT; digit3<=TWO; end
      16'd2870: begin digit0<=ZERO; digit1<=SEVEN; digit2<=EIGHT; digit3<=TWO; end
      16'd2871: begin digit0<=ONE; digit1<=SEVEN; digit2<=EIGHT; digit3<=TWO; end
      16'd2872: begin digit0<=TWO; digit1<=SEVEN; digit2<=EIGHT; digit3<=TWO; end
      16'd2873: begin digit0<=THREE; digit1<=SEVEN; digit2<=EIGHT; digit3<=TWO; end
      16'd2874: begin digit0<=FOUR; digit1<=SEVEN; digit2<=EIGHT; digit3<=TWO; end
      16'd2875: begin digit0<=FIVE; digit1<=SEVEN; digit2<=EIGHT; digit3<=TWO; end
      16'd2876: begin digit0<=SIX; digit1<=SEVEN; digit2<=EIGHT; digit3<=TWO; end
      16'd2877: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=EIGHT; digit3<=TWO; end
      16'd2878: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=EIGHT; digit3<=TWO; end
      16'd2879: begin digit0<=NINE; digit1<=SEVEN; digit2<=EIGHT; digit3<=TWO; end
      16'd2880: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=TWO; end
      16'd2881: begin digit0<=ONE; digit1<=EIGHT; digit2<=EIGHT; digit3<=TWO; end
      16'd2882: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=TWO; end
      16'd2883: begin digit0<=THREE; digit1<=EIGHT; digit2<=EIGHT; digit3<=TWO; end
      16'd2884: begin digit0<=FOUR; digit1<=EIGHT; digit2<=EIGHT; digit3<=TWO; end
      16'd2885: begin digit0<=FIVE; digit1<=EIGHT; digit2<=EIGHT; digit3<=TWO; end
      16'd2886: begin digit0<=SIX; digit1<=EIGHT; digit2<=EIGHT; digit3<=TWO; end
      16'd2887: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=EIGHT; digit3<=TWO; end
      16'd2888: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=EIGHT; digit3<=TWO; end
      16'd2889: begin digit0<=NINE; digit1<=EIGHT; digit2<=EIGHT; digit3<=TWO; end
      16'd2890: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=TWO; end
      16'd2891: begin digit0<=ONE; digit1<=NINE; digit2<=EIGHT; digit3<=TWO; end
      16'd2892: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=TWO; end
      16'd2893: begin digit0<=THREE; digit1<=NINE; digit2<=EIGHT; digit3<=TWO; end
      16'd2894: begin digit0<=FOUR; digit1<=NINE; digit2<=EIGHT; digit3<=TWO; end
      16'd2895: begin digit0<=FIVE; digit1<=NINE; digit2<=EIGHT; digit3<=TWO; end
      16'd2896: begin digit0<=SIX; digit1<=NINE; digit2<=EIGHT; digit3<=TWO; end
      16'd2897: begin digit0<=SEVEN; digit1<=NINE; digit2<=EIGHT; digit3<=TWO; end
      16'd2898: begin digit0<=EIGHT; digit1<=NINE; digit2<=EIGHT; digit3<=TWO; end
      16'd2899: begin digit0<=NINE; digit1<=NINE; digit2<=EIGHT; digit3<=TWO; end
	  16'd2900: begin digit0<=ZERO; digit1<=ZERO; digit2<=NINE; digit3<=TWO; end
      16'd2901: begin digit0<=ONE; digit1<=ZERO; digit2<=NINE; digit3<=TWO; end
      16'd2902: begin digit0<=TWO; digit1<=ZERO; digit2<=NINE; digit3<=TWO; end
      16'd2903: begin digit0<=THREE; digit1<=ZERO; digit2<=NINE; digit3<=TWO; end
      16'd2904: begin digit0<=FOUR; digit1<=ZERO; digit2<=NINE; digit3<=TWO; end
      16'd2905: begin digit0<=FIVE; digit1<=ZERO; digit2<=NINE; digit3<=TWO; end
      16'd2906: begin digit0<=SIX; digit1<=ZERO; digit2<=NINE; digit3<=TWO; end
      16'd2907: begin digit0<=SEVEN; digit1<=ZERO; digit2<=NINE; digit3<=TWO; end
      16'd2908: begin digit0<=EIGHT; digit1<=ZERO; digit2<=NINE; digit3<=TWO; end
      16'd2909: begin digit0<=NINE; digit1<=ZERO; digit2<=NINE; digit3<=TWO; end
      16'd2910: begin digit0<=ZERO; digit1<=ONE; digit2<=NINE; digit3<=TWO; end
      16'd2911: begin digit0<=ONE; digit1<=ONE; digit2<=NINE; digit3<=TWO; end
      16'd2912: begin digit0<=TWO; digit1<=ONE; digit2<=NINE; digit3<=TWO; end
      16'd2913: begin digit0<=THREE; digit1<=ONE; digit2<=NINE; digit3<=TWO; end
      16'd2914: begin digit0<=FOUR; digit1<=ONE; digit2<=NINE; digit3<=TWO; end
      16'd2915: begin digit0<=FIVE; digit1<=ONE; digit2<=NINE; digit3<=TWO; end
      16'd2916: begin digit0<=SIX; digit1<=ONE; digit2<=NINE; digit3<=TWO; end
      16'd2917: begin digit0<=SEVEN; digit1<=ONE; digit2<=NINE; digit3<=TWO; end
      16'd2918: begin digit0<=EIGHT; digit1<=ONE; digit2<=NINE; digit3<=TWO; end
      16'd2919: begin digit0<=NINE; digit1<=ONE; digit2<=NINE; digit3<=TWO; end
      16'd2920: begin digit0<=ZERO; digit1<=TWO; digit2<=NINE; digit3<=TWO; end
      16'd2921: begin digit0<=ONE; digit1<=TWO; digit2<=NINE; digit3<=TWO; end
      16'd2922: begin digit0<=TWO; digit1<=TWO; digit2<=NINE; digit3<=TWO; end
      16'd2923: begin digit0<=THREE; digit1<=TWO; digit2<=NINE; digit3<=TWO; end
      16'd2924: begin digit0<=FOUR; digit1<=TWO; digit2<=NINE; digit3<=TWO; end
      16'd2925: begin digit0<=FIVE; digit1<=TWO; digit2<=NINE; digit3<=TWO; end
      16'd2926: begin digit0<=SIX; digit1<=TWO; digit2<=NINE; digit3<=TWO; end
      16'd2927: begin digit0<=SEVEN; digit1<=TWO; digit2<=NINE; digit3<=TWO; end
      16'd2928: begin digit0<=EIGHT; digit1<=TWO; digit2<=NINE; digit3<=TWO; end
      16'd2929: begin digit0<=NINE; digit1<=TWO; digit2<=NINE; digit3<=TWO; end
      16'd2930: begin digit0<=ZERO; digit1<=THREE; digit2<=NINE; digit3<=TWO; end
      16'd2931: begin digit0<=ONE; digit1<=THREE; digit2<=NINE; digit3<=TWO; end
      16'd2932: begin digit0<=TWO; digit1<=THREE; digit2<=NINE; digit3<=TWO; end
      16'd2933: begin digit0<=THREE; digit1<=THREE; digit2<=NINE; digit3<=TWO; end
      16'd2934: begin digit0<=FOUR; digit1<=THREE; digit2<=NINE; digit3<=TWO; end
      16'd2935: begin digit0<=FIVE; digit1<=THREE; digit2<=NINE; digit3<=TWO; end
      16'd2936: begin digit0<=SIX; digit1<=THREE; digit2<=NINE; digit3<=TWO; end
      16'd2937: begin digit0<=SEVEN; digit1<=THREE; digit2<=NINE; digit3<=TWO; end
      16'd2938: begin digit0<=EIGHT; digit1<=THREE; digit2<=NINE; digit3<=TWO; end
      16'd2939: begin digit0<=NINE; digit1<=THREE; digit2<=NINE; digit3<=TWO; end
      16'd2940: begin digit0<=ZERO; digit1<=FOUR; digit2<=NINE; digit3<=TWO; end
      16'd2941: begin digit0<=ONE; digit1<=FOUR; digit2<=NINE; digit3<=TWO; end
      16'd2942: begin digit0<=TWO; digit1<=FOUR; digit2<=NINE; digit3<=TWO; end
      16'd2943: begin digit0<=THREE; digit1<=FOUR; digit2<=NINE; digit3<=TWO; end
      16'd2944: begin digit0<=FOUR; digit1<=FOUR; digit2<=NINE; digit3<=TWO; end
      16'd2945: begin digit0<=FIVE; digit1<=FOUR; digit2<=NINE; digit3<=TWO; end
      16'd2946: begin digit0<=SIX; digit1<=FOUR; digit2<=NINE; digit3<=TWO; end
      16'd2947: begin digit0<=SEVEN; digit1<=FOUR; digit2<=NINE; digit3<=TWO; end
      16'd2948: begin digit0<=EIGHT; digit1<=FOUR; digit2<=NINE; digit3<=TWO; end
      16'd2949: begin digit0<=NINE; digit1<=FOUR; digit2<=NINE; digit3<=TWO; end
      16'd2950: begin digit0<=ZERO; digit1<=FIVE; digit2<=NINE; digit3<=TWO; end
      16'd2951: begin digit0<=ONE; digit1<=FIVE; digit2<=NINE; digit3<=TWO; end
      16'd2952: begin digit0<=TWO; digit1<=FIVE; digit2<=NINE; digit3<=TWO; end
      16'd2953: begin digit0<=THREE; digit1<=FIVE; digit2<=NINE; digit3<=TWO; end
      16'd2954: begin digit0<=FOUR; digit1<=FIVE; digit2<=NINE; digit3<=TWO; end
      16'd2955: begin digit0<=FIVE; digit1<=FIVE; digit2<=NINE; digit3<=TWO; end
      16'd2956: begin digit0<=SIX; digit1<=FIVE; digit2<=NINE; digit3<=TWO; end
      16'd2957: begin digit0<=SEVEN; digit1<=FIVE; digit2<=NINE; digit3<=TWO; end
      16'd2958: begin digit0<=EIGHT; digit1<=FIVE; digit2<=NINE; digit3<=TWO; end
      16'd2959: begin digit0<=NINE; digit1<=FIVE; digit2<=NINE; digit3<=TWO; end
      16'd2960: begin digit0<=ZERO; digit1<=SIX; digit2<=NINE; digit3<=TWO; end
      16'd2961: begin digit0<=ONE; digit1<=SIX; digit2<=NINE; digit3<=TWO; end
      16'd2962: begin digit0<=TWO; digit1<=SIX; digit2<=NINE; digit3<=TWO; end
      16'd2963: begin digit0<=THREE; digit1<=SIX; digit2<=NINE; digit3<=TWO; end
      16'd2964: begin digit0<=FOUR; digit1<=SIX; digit2<=NINE; digit3<=TWO; end
      16'd2965: begin digit0<=FIVE; digit1<=SIX; digit2<=NINE; digit3<=TWO; end
      16'd2966: begin digit0<=SIX; digit1<=SIX; digit2<=NINE; digit3<=TWO; end
      16'd2967: begin digit0<=SEVEN; digit1<=SIX; digit2<=NINE; digit3<=TWO; end
      16'd2968: begin digit0<=EIGHT; digit1<=SIX; digit2<=NINE; digit3<=TWO; end
      16'd2969: begin digit0<=NINE; digit1<=SIX; digit2<=NINE; digit3<=TWO; end
      16'd2970: begin digit0<=ZERO; digit1<=SEVEN; digit2<=NINE; digit3<=TWO; end
      16'd2971: begin digit0<=ONE; digit1<=SEVEN; digit2<=NINE; digit3<=TWO; end
      16'd2972: begin digit0<=TWO; digit1<=SEVEN; digit2<=NINE; digit3<=TWO; end
      16'd2973: begin digit0<=THREE; digit1<=SEVEN; digit2<=NINE; digit3<=TWO; end
      16'd2974: begin digit0<=FOUR; digit1<=SEVEN; digit2<=NINE; digit3<=TWO; end
      16'd2975: begin digit0<=FIVE; digit1<=SEVEN; digit2<=NINE; digit3<=TWO; end
      16'd2976: begin digit0<=SIX; digit1<=SEVEN; digit2<=NINE; digit3<=TWO; end
      16'd2977: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=NINE; digit3<=TWO; end
      16'd2978: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=NINE; digit3<=TWO; end
      16'd2979: begin digit0<=NINE; digit1<=SEVEN; digit2<=NINE; digit3<=TWO; end
      16'd2980: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=TWO; end
      16'd2981: begin digit0<=ONE; digit1<=EIGHT; digit2<=NINE; digit3<=TWO; end
      16'd2982: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=TWO; end
      16'd2983: begin digit0<=THREE; digit1<=EIGHT; digit2<=NINE; digit3<=TWO; end
      16'd2984: begin digit0<=FOUR; digit1<=EIGHT; digit2<=NINE; digit3<=TWO; end
      16'd2985: begin digit0<=FIVE; digit1<=EIGHT; digit2<=NINE; digit3<=TWO; end
      16'd2986: begin digit0<=SIX; digit1<=EIGHT; digit2<=NINE; digit3<=TWO; end
      16'd2987: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=NINE; digit3<=TWO; end
      16'd2988: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=NINE; digit3<=TWO; end
      16'd2989: begin digit0<=NINE; digit1<=EIGHT; digit2<=NINE; digit3<=TWO; end
      16'd2990: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=TWO; end
      16'd2991: begin digit0<=ONE; digit1<=NINE; digit2<=NINE; digit3<=TWO; end
      16'd2992: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=TWO; end
      16'd2993: begin digit0<=THREE; digit1<=NINE; digit2<=NINE; digit3<=TWO; end
      16'd2994: begin digit0<=FOUR; digit1<=NINE; digit2<=NINE; digit3<=TWO; end
      16'd2995: begin digit0<=FIVE; digit1<=NINE; digit2<=NINE; digit3<=TWO; end
      16'd2996: begin digit0<=SIX; digit1<=NINE; digit2<=NINE; digit3<=TWO; end
      16'd2997: begin digit0<=SEVEN; digit1<=NINE; digit2<=NINE; digit3<=TWO; end
      16'd2998: begin digit0<=EIGHT; digit1<=NINE; digit2<=NINE; digit3<=TWO; end
      16'd2999: begin digit0<=NINE; digit1<=NINE; digit2<=NINE; digit3<=TWO; end
	  16'd3000: begin digit0<=ZERO; digit1<=ZERO; digit2<=ZERO; digit3<=THREE; end
      16'd3001: begin digit0<=ONE; digit1<=ZERO; digit2<=ZERO; digit3<=THREE; end
      16'd3002: begin digit0<=TWO; digit1<=ZERO; digit2<=ZERO; digit3<=THREE; end
      16'd3003: begin digit0<=THREE; digit1<=ZERO; digit2<=ZERO; digit3<=THREE; end
      16'd3004: begin digit0<=FOUR; digit1<=ZERO; digit2<=ZERO; digit3<=THREE; end
      16'd3005: begin digit0<=FIVE; digit1<=ZERO; digit2<=ZERO; digit3<=THREE; end
      16'd3006: begin digit0<=SIX; digit1<=ZERO; digit2<=ZERO; digit3<=THREE; end
      16'd3007: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ZERO; digit3<=THREE; end
      16'd3008: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ZERO; digit3<=THREE; end
      16'd3009: begin digit0<=NINE; digit1<=ZERO; digit2<=ZERO; digit3<=THREE; end
      16'd3010: begin digit0<=ZERO; digit1<=ONE; digit2<=ZERO; digit3<=THREE; end
      16'd3011: begin digit0<=ONE; digit1<=ONE; digit2<=ZERO; digit3<=THREE; end
      16'd3012: begin digit0<=TWO; digit1<=ONE; digit2<=ZERO; digit3<=THREE; end
      16'd3013: begin digit0<=THREE; digit1<=ONE; digit2<=ZERO; digit3<=THREE; end
      16'd3014: begin digit0<=FOUR; digit1<=ONE; digit2<=ZERO; digit3<=THREE; end
      16'd3015: begin digit0<=FIVE; digit1<=ONE; digit2<=ZERO; digit3<=THREE; end
      16'd3016: begin digit0<=SIX; digit1<=ONE; digit2<=ZERO; digit3<=THREE; end
      16'd3017: begin digit0<=SEVEN; digit1<=ONE; digit2<=ZERO; digit3<=THREE; end
      16'd3018: begin digit0<=EIGHT; digit1<=ONE; digit2<=ZERO; digit3<=THREE; end
      16'd3019: begin digit0<=NINE; digit1<=ONE; digit2<=ZERO; digit3<=THREE; end
      16'd3020: begin digit0<=ZERO; digit1<=TWO; digit2<=ZERO; digit3<=THREE; end
      16'd3021: begin digit0<=ONE; digit1<=TWO; digit2<=ZERO; digit3<=THREE; end
      16'd3022: begin digit0<=TWO; digit1<=TWO; digit2<=ZERO; digit3<=THREE; end
      16'd3023: begin digit0<=THREE; digit1<=TWO; digit2<=ZERO; digit3<=THREE; end
      16'd3024: begin digit0<=FOUR; digit1<=TWO; digit2<=ZERO; digit3<=THREE; end
      16'd3025: begin digit0<=FIVE; digit1<=TWO; digit2<=ZERO; digit3<=THREE; end
      16'd3026: begin digit0<=SIX; digit1<=TWO; digit2<=ZERO; digit3<=THREE; end
      16'd3027: begin digit0<=SEVEN; digit1<=TWO; digit2<=ZERO; digit3<=THREE; end
      16'd3028: begin digit0<=EIGHT; digit1<=TWO; digit2<=ZERO; digit3<=THREE; end
      16'd3029: begin digit0<=NINE; digit1<=TWO; digit2<=ZERO; digit3<=THREE; end
      16'd3030: begin digit0<=ZERO; digit1<=THREE; digit2<=ZERO; digit3<=THREE; end
      16'd3031: begin digit0<=ONE; digit1<=THREE; digit2<=ZERO; digit3<=THREE; end
      16'd3032: begin digit0<=TWO; digit1<=THREE; digit2<=ZERO; digit3<=THREE; end
      16'd3033: begin digit0<=THREE; digit1<=THREE; digit2<=ZERO; digit3<=THREE; end
      16'd3034: begin digit0<=FOUR; digit1<=THREE; digit2<=ZERO; digit3<=THREE; end
      16'd3035: begin digit0<=FIVE; digit1<=THREE; digit2<=ZERO; digit3<=THREE; end
      16'd3036: begin digit0<=SIX; digit1<=THREE; digit2<=ZERO; digit3<=THREE; end
      16'd3037: begin digit0<=SEVEN; digit1<=THREE; digit2<=ZERO; digit3<=THREE; end
      16'd3038: begin digit0<=EIGHT; digit1<=THREE; digit2<=ZERO; digit3<=THREE; end
      16'd3039: begin digit0<=NINE; digit1<=THREE; digit2<=ZERO; digit3<=THREE; end
      16'd3040: begin digit0<=ZERO; digit1<=FOUR; digit2<=ZERO; digit3<=THREE; end
      16'd3041: begin digit0<=ONE; digit1<=FOUR; digit2<=ZERO; digit3<=THREE; end
      16'd3042: begin digit0<=TWO; digit1<=FOUR; digit2<=ZERO; digit3<=THREE; end
      16'd3043: begin digit0<=THREE; digit1<=FOUR; digit2<=ZERO; digit3<=THREE; end
      16'd3044: begin digit0<=FOUR; digit1<=FOUR; digit2<=ZERO; digit3<=THREE; end
      16'd3045: begin digit0<=FIVE; digit1<=FOUR; digit2<=ZERO; digit3<=THREE; end
      16'd3046: begin digit0<=SIX; digit1<=FOUR; digit2<=ZERO; digit3<=THREE; end
      16'd3047: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ZERO; digit3<=THREE; end
      16'd3048: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ZERO; digit3<=THREE; end
      16'd3049: begin digit0<=NINE; digit1<=FOUR; digit2<=ZERO; digit3<=THREE; end
      16'd3050: begin digit0<=ZERO; digit1<=FIVE; digit2<=ZERO; digit3<=THREE; end
      16'd3051: begin digit0<=ONE; digit1<=FIVE; digit2<=ZERO; digit3<=THREE; end
      16'd3052: begin digit0<=TWO; digit1<=FIVE; digit2<=ZERO; digit3<=THREE; end
      16'd3053: begin digit0<=THREE; digit1<=FIVE; digit2<=ZERO; digit3<=THREE; end
      16'd3054: begin digit0<=FOUR; digit1<=FIVE; digit2<=ZERO; digit3<=THREE; end
      16'd3055: begin digit0<=FIVE; digit1<=FIVE; digit2<=ZERO; digit3<=THREE; end
      16'd3056: begin digit0<=SIX; digit1<=FIVE; digit2<=ZERO; digit3<=THREE; end
      16'd3057: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ZERO; digit3<=THREE; end
      16'd3058: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ZERO; digit3<=THREE; end
      16'd3059: begin digit0<=NINE; digit1<=FIVE; digit2<=ZERO; digit3<=THREE; end
      16'd3060: begin digit0<=ZERO; digit1<=SIX; digit2<=ZERO; digit3<=THREE; end
      16'd3061: begin digit0<=ONE; digit1<=SIX; digit2<=ZERO; digit3<=THREE; end
      16'd3062: begin digit0<=TWO; digit1<=SIX; digit2<=ZERO; digit3<=THREE; end
      16'd3063: begin digit0<=THREE; digit1<=SIX; digit2<=ZERO; digit3<=THREE; end
      16'd3064: begin digit0<=FOUR; digit1<=SIX; digit2<=ZERO; digit3<=THREE; end
      16'd3065: begin digit0<=FIVE; digit1<=SIX; digit2<=ZERO; digit3<=THREE; end
      16'd3066: begin digit0<=SIX; digit1<=SIX; digit2<=ZERO; digit3<=THREE; end
      16'd3067: begin digit0<=SEVEN; digit1<=SIX; digit2<=ZERO; digit3<=THREE; end
      16'd3068: begin digit0<=EIGHT; digit1<=SIX; digit2<=ZERO; digit3<=THREE; end
      16'd3069: begin digit0<=NINE; digit1<=SIX; digit2<=ZERO; digit3<=THREE; end
      16'd3070: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ZERO; digit3<=THREE; end
      16'd3071: begin digit0<=ONE; digit1<=SEVEN; digit2<=ZERO; digit3<=THREE; end
      16'd3072: begin digit0<=TWO; digit1<=SEVEN; digit2<=ZERO; digit3<=THREE; end
      16'd3073: begin digit0<=THREE; digit1<=SEVEN; digit2<=ZERO; digit3<=THREE; end
      16'd3074: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ZERO; digit3<=THREE; end
      16'd3075: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ZERO; digit3<=THREE; end
      16'd3076: begin digit0<=SIX; digit1<=SEVEN; digit2<=ZERO; digit3<=THREE; end
      16'd3077: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ZERO; digit3<=THREE; end
      16'd3078: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ZERO; digit3<=THREE; end
      16'd3079: begin digit0<=NINE; digit1<=SEVEN; digit2<=ZERO; digit3<=THREE; end
      16'd3080: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ZERO; digit3<=THREE; end
      16'd3081: begin digit0<=ONE; digit1<=EIGHT; digit2<=ZERO; digit3<=THREE; end
      16'd3082: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ZERO; digit3<=THREE; end
      16'd3083: begin digit0<=THREE; digit1<=EIGHT; digit2<=ZERO; digit3<=THREE; end
      16'd3084: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ZERO; digit3<=THREE; end
      16'd3085: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ZERO; digit3<=THREE; end
      16'd3086: begin digit0<=SIX; digit1<=EIGHT; digit2<=ZERO; digit3<=THREE; end
      16'd3087: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ZERO; digit3<=THREE; end
      16'd3088: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ZERO; digit3<=THREE; end
      16'd3089: begin digit0<=NINE; digit1<=EIGHT; digit2<=ZERO; digit3<=THREE; end
      16'd3090: begin digit0<=ZERO; digit1<=NINE; digit2<=ZERO; digit3<=THREE; end
      16'd3091: begin digit0<=ONE; digit1<=NINE; digit2<=ZERO; digit3<=THREE; end
      16'd3092: begin digit0<=ZERO; digit1<=NINE; digit2<=ZERO; digit3<=THREE; end
      16'd3093: begin digit0<=THREE; digit1<=NINE; digit2<=ZERO; digit3<=THREE; end
      16'd3094: begin digit0<=FOUR; digit1<=NINE; digit2<=ZERO; digit3<=THREE; end
      16'd3095: begin digit0<=FIVE; digit1<=NINE; digit2<=ZERO; digit3<=THREE; end
      16'd3096: begin digit0<=SIX; digit1<=NINE; digit2<=ZERO; digit3<=THREE; end
      16'd3097: begin digit0<=SEVEN; digit1<=NINE; digit2<=ZERO; digit3<=THREE; end
      16'd3098: begin digit0<=EIGHT; digit1<=NINE; digit2<=ZERO; digit3<=THREE; end
      16'd3099: begin digit0<=NINE; digit1<=NINE; digit2<=ZERO; digit3<=THREE; end
	  16'd3100: begin digit0<=ZERO; digit1<=ZERO; digit2<=ONE; digit3<=THREE; end
      16'd3101: begin digit0<=ONE; digit1<=ZERO; digit2<=ONE; digit3<=THREE; end
      16'd3102: begin digit0<=TWO; digit1<=ZERO; digit2<=ONE; digit3<=THREE; end
      16'd3103: begin digit0<=THREE; digit1<=ZERO; digit2<=ONE; digit3<=THREE; end
      16'd3104: begin digit0<=FOUR; digit1<=ZERO; digit2<=ONE; digit3<=THREE; end
      16'd3105: begin digit0<=FIVE; digit1<=ZERO; digit2<=ONE; digit3<=THREE; end
      16'd3106: begin digit0<=SIX; digit1<=ZERO; digit2<=ONE; digit3<=THREE; end
      16'd3107: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ONE; digit3<=THREE; end
      16'd3108: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ONE; digit3<=THREE; end
      16'd3109: begin digit0<=NINE; digit1<=ZERO; digit2<=ONE; digit3<=THREE; end
      16'd3110: begin digit0<=ZERO; digit1<=ONE; digit2<=ONE; digit3<=THREE; end
      16'd3111: begin digit0<=ONE; digit1<=ONE; digit2<=ONE; digit3<=THREE; end
      16'd3112: begin digit0<=TWO; digit1<=ONE; digit2<=ONE; digit3<=THREE; end
      16'd3113: begin digit0<=THREE; digit1<=ONE; digit2<=ONE; digit3<=THREE; end
      16'd3114: begin digit0<=FOUR; digit1<=ONE; digit2<=ONE; digit3<=THREE; end
      16'd3115: begin digit0<=FIVE; digit1<=ONE; digit2<=ONE; digit3<=THREE; end
      16'd3116: begin digit0<=SIX; digit1<=ONE; digit2<=ONE; digit3<=THREE; end
      16'd3117: begin digit0<=SEVEN; digit1<=ONE; digit2<=ONE; digit3<=THREE; end
      16'd3118: begin digit0<=EIGHT; digit1<=ONE; digit2<=ONE; digit3<=THREE; end
      16'd3119: begin digit0<=NINE; digit1<=ONE; digit2<=ONE; digit3<=THREE; end
      16'd3120: begin digit0<=ZERO; digit1<=TWO; digit2<=ONE; digit3<=THREE; end
      16'd3121: begin digit0<=ONE; digit1<=TWO; digit2<=ONE; digit3<=THREE; end
      16'd3122: begin digit0<=TWO; digit1<=TWO; digit2<=ONE; digit3<=THREE; end
      16'd3123: begin digit0<=THREE; digit1<=TWO; digit2<=ONE; digit3<=THREE; end
      16'd3124: begin digit0<=FOUR; digit1<=TWO; digit2<=ONE; digit3<=THREE; end
      16'd3125: begin digit0<=FIVE; digit1<=TWO; digit2<=ONE; digit3<=THREE; end
      16'd3126: begin digit0<=SIX; digit1<=TWO; digit2<=ONE; digit3<=THREE; end
      16'd3127: begin digit0<=SEVEN; digit1<=TWO; digit2<=ONE; digit3<=THREE; end
      16'd3128: begin digit0<=EIGHT; digit1<=TWO; digit2<=ONE; digit3<=THREE; end
      16'd3129: begin digit0<=NINE; digit1<=TWO; digit2<=ONE; digit3<=THREE; end
      16'd3130: begin digit0<=ZERO; digit1<=THREE; digit2<=ONE; digit3<=THREE; end
      16'd3131: begin digit0<=ONE; digit1<=THREE; digit2<=ONE; digit3<=THREE; end
      16'd3132: begin digit0<=TWO; digit1<=THREE; digit2<=ONE; digit3<=THREE; end
      16'd3133: begin digit0<=THREE; digit1<=THREE; digit2<=ONE; digit3<=THREE; end
      16'd3134: begin digit0<=FOUR; digit1<=THREE; digit2<=ONE; digit3<=THREE; end
      16'd3135: begin digit0<=FIVE; digit1<=THREE; digit2<=ONE; digit3<=THREE; end
      16'd3136: begin digit0<=SIX; digit1<=THREE; digit2<=ONE; digit3<=THREE; end
      16'd3137: begin digit0<=SEVEN; digit1<=THREE; digit2<=ONE; digit3<=THREE; end
      16'd3138: begin digit0<=EIGHT; digit1<=THREE; digit2<=ONE; digit3<=THREE; end
      16'd3139: begin digit0<=NINE; digit1<=THREE; digit2<=ONE; digit3<=THREE; end
      16'd3140: begin digit0<=ZERO; digit1<=FOUR; digit2<=ONE; digit3<=THREE; end
      16'd3141: begin digit0<=ONE; digit1<=FOUR; digit2<=ONE; digit3<=THREE; end
      16'd3142: begin digit0<=TWO; digit1<=FOUR; digit2<=ONE; digit3<=THREE; end
      16'd3143: begin digit0<=THREE; digit1<=FOUR; digit2<=ONE; digit3<=THREE; end
      16'd3144: begin digit0<=FOUR; digit1<=FOUR; digit2<=ONE; digit3<=THREE; end
      16'd3145: begin digit0<=FIVE; digit1<=FOUR; digit2<=ONE; digit3<=THREE; end
      16'd3146: begin digit0<=SIX; digit1<=FOUR; digit2<=ONE; digit3<=THREE; end
      16'd3147: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ONE; digit3<=THREE; end
      16'd3148: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ONE; digit3<=THREE; end
      16'd3149: begin digit0<=NINE; digit1<=FOUR; digit2<=ONE; digit3<=THREE; end
      16'd3150: begin digit0<=ZERO; digit1<=FIVE; digit2<=ONE; digit3<=THREE; end
      16'd3151: begin digit0<=ONE; digit1<=FIVE; digit2<=ONE; digit3<=THREE; end
      16'd3152: begin digit0<=TWO; digit1<=FIVE; digit2<=ONE; digit3<=THREE; end
      16'd3153: begin digit0<=THREE; digit1<=FIVE; digit2<=ONE; digit3<=THREE; end
      16'd3154: begin digit0<=FOUR; digit1<=FIVE; digit2<=ONE; digit3<=THREE; end
      16'd3155: begin digit0<=FIVE; digit1<=FIVE; digit2<=ONE; digit3<=THREE; end
      16'd3156: begin digit0<=SIX; digit1<=FIVE; digit2<=ONE; digit3<=THREE; end
      16'd3157: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ONE; digit3<=THREE; end
      16'd3158: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ONE; digit3<=THREE; end
      16'd3159: begin digit0<=NINE; digit1<=FIVE; digit2<=ONE; digit3<=THREE; end
      16'd3160: begin digit0<=ZERO; digit1<=SIX; digit2<=ONE; digit3<=THREE; end
      16'd3161: begin digit0<=ONE; digit1<=SIX; digit2<=ONE; digit3<=THREE; end
      16'd3162: begin digit0<=TWO; digit1<=SIX; digit2<=ONE; digit3<=THREE; end
      16'd3163: begin digit0<=THREE; digit1<=SIX; digit2<=ONE; digit3<=THREE; end
      16'd3164: begin digit0<=FOUR; digit1<=SIX; digit2<=ONE; digit3<=THREE; end
      16'd3165: begin digit0<=FIVE; digit1<=SIX; digit2<=ONE; digit3<=THREE; end
      16'd3166: begin digit0<=SIX; digit1<=SIX; digit2<=ONE; digit3<=THREE; end
      16'd3167: begin digit0<=SEVEN; digit1<=SIX; digit2<=ONE; digit3<=THREE; end
      16'd3168: begin digit0<=EIGHT; digit1<=SIX; digit2<=ONE; digit3<=THREE; end
      16'd3169: begin digit0<=NINE; digit1<=SIX; digit2<=ONE; digit3<=THREE; end
      16'd3170: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ONE; digit3<=THREE; end
      16'd3171: begin digit0<=ONE; digit1<=SEVEN; digit2<=ONE; digit3<=THREE; end
      16'd3172: begin digit0<=TWO; digit1<=SEVEN; digit2<=ONE; digit3<=THREE; end
      16'd3173: begin digit0<=THREE; digit1<=SEVEN; digit2<=ONE; digit3<=THREE; end
      16'd3174: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ONE; digit3<=THREE; end
      16'd3175: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ONE; digit3<=THREE; end
      16'd3176: begin digit0<=SIX; digit1<=SEVEN; digit2<=ONE; digit3<=THREE; end
      16'd3177: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ONE; digit3<=THREE; end
      16'd3178: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ONE; digit3<=THREE; end
      16'd3179: begin digit0<=NINE; digit1<=SEVEN; digit2<=ONE; digit3<=THREE; end
      16'd3180: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=THREE; end
      16'd3181: begin digit0<=ONE; digit1<=EIGHT; digit2<=ONE; digit3<=THREE; end
      16'd3182: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=THREE; end
      16'd3183: begin digit0<=THREE; digit1<=EIGHT; digit2<=ONE; digit3<=THREE; end
      16'd3184: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ONE; digit3<=THREE; end
      16'd3185: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ONE; digit3<=THREE; end
      16'd3186: begin digit0<=SIX; digit1<=EIGHT; digit2<=ONE; digit3<=THREE; end
      16'd3187: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ONE; digit3<=THREE; end
      16'd3188: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ONE; digit3<=THREE; end
      16'd3189: begin digit0<=NINE; digit1<=EIGHT; digit2<=ONE; digit3<=THREE; end
      16'd3190: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=THREE; end
      16'd3191: begin digit0<=ONE; digit1<=NINE; digit2<=ONE; digit3<=THREE; end
      16'd3192: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=THREE; end
      16'd3193: begin digit0<=THREE; digit1<=NINE; digit2<=ONE; digit3<=THREE; end
      16'd3194: begin digit0<=FOUR; digit1<=NINE; digit2<=ONE; digit3<=THREE; end
      16'd3195: begin digit0<=FIVE; digit1<=NINE; digit2<=ONE; digit3<=THREE; end
      16'd3196: begin digit0<=SIX; digit1<=NINE; digit2<=ONE; digit3<=THREE; end
      16'd3197: begin digit0<=SEVEN; digit1<=NINE; digit2<=ONE; digit3<=THREE; end
      16'd3198: begin digit0<=EIGHT; digit1<=NINE; digit2<=ONE; digit3<=THREE; end
      16'd3199: begin digit0<=NINE; digit1<=NINE; digit2<=ONE; digit3<=THREE; end
	  16'd3200: begin digit0<=ZERO; digit1<=ZERO; digit2<=TWO; digit3<=THREE; end
      16'd3201: begin digit0<=ONE; digit1<=ZERO; digit2<=TWO; digit3<=THREE; end
      16'd3202: begin digit0<=TWO; digit1<=ZERO; digit2<=TWO; digit3<=THREE; end
      16'd3203: begin digit0<=THREE; digit1<=ZERO; digit2<=TWO; digit3<=THREE; end
      16'd3204: begin digit0<=FOUR; digit1<=ZERO; digit2<=TWO; digit3<=THREE; end
      16'd3205: begin digit0<=FIVE; digit1<=ZERO; digit2<=TWO; digit3<=THREE; end
      16'd3206: begin digit0<=SIX; digit1<=ZERO; digit2<=TWO; digit3<=THREE; end
      16'd3207: begin digit0<=SEVEN; digit1<=ZERO; digit2<=TWO; digit3<=THREE; end
      16'd3208: begin digit0<=EIGHT; digit1<=ZERO; digit2<=TWO; digit3<=THREE; end
      16'd3209: begin digit0<=NINE; digit1<=ZERO; digit2<=TWO; digit3<=THREE; end
      16'd3210: begin digit0<=ZERO; digit1<=ONE; digit2<=TWO; digit3<=THREE; end
      16'd3211: begin digit0<=ONE; digit1<=ONE; digit2<=TWO; digit3<=THREE; end
      16'd3212: begin digit0<=TWO; digit1<=ONE; digit2<=TWO; digit3<=THREE; end
      16'd3213: begin digit0<=THREE; digit1<=ONE; digit2<=TWO; digit3<=THREE; end
      16'd3214: begin digit0<=FOUR; digit1<=ONE; digit2<=TWO; digit3<=THREE; end
      16'd3215: begin digit0<=FIVE; digit1<=ONE; digit2<=TWO; digit3<=THREE; end
      16'd3216: begin digit0<=SIX; digit1<=ONE; digit2<=TWO; digit3<=THREE; end
      16'd3217: begin digit0<=SEVEN; digit1<=ONE; digit2<=TWO; digit3<=THREE; end
      16'd3218: begin digit0<=EIGHT; digit1<=ONE; digit2<=TWO; digit3<=THREE; end
      16'd3219: begin digit0<=NINE; digit1<=ONE; digit2<=TWO; digit3<=THREE; end
      16'd3220: begin digit0<=ZERO; digit1<=TWO; digit2<=TWO; digit3<=THREE; end
      16'd3221: begin digit0<=ONE; digit1<=TWO; digit2<=TWO; digit3<=THREE; end
      16'd3222: begin digit0<=TWO; digit1<=TWO; digit2<=TWO; digit3<=THREE; end
      16'd3223: begin digit0<=THREE; digit1<=TWO; digit2<=TWO; digit3<=THREE; end
      16'd3224: begin digit0<=FOUR; digit1<=TWO; digit2<=TWO; digit3<=THREE; end
      16'd3225: begin digit0<=FIVE; digit1<=TWO; digit2<=TWO; digit3<=THREE; end
      16'd3226: begin digit0<=SIX; digit1<=TWO; digit2<=TWO; digit3<=THREE; end
      16'd3227: begin digit0<=SEVEN; digit1<=TWO; digit2<=TWO; digit3<=THREE; end
      16'd3228: begin digit0<=EIGHT; digit1<=TWO; digit2<=TWO; digit3<=THREE; end
      16'd3229: begin digit0<=NINE; digit1<=TWO; digit2<=TWO; digit3<=THREE; end
      16'd3230: begin digit0<=ZERO; digit1<=THREE; digit2<=TWO; digit3<=THREE; end
      16'd3231: begin digit0<=ONE; digit1<=THREE; digit2<=TWO; digit3<=THREE; end
      16'd3232: begin digit0<=TWO; digit1<=THREE; digit2<=TWO; digit3<=THREE; end
      16'd3233: begin digit0<=THREE; digit1<=THREE; digit2<=TWO; digit3<=THREE; end
      16'd3234: begin digit0<=FOUR; digit1<=THREE; digit2<=TWO; digit3<=THREE; end
      16'd3235: begin digit0<=FIVE; digit1<=THREE; digit2<=TWO; digit3<=THREE; end
      16'd3236: begin digit0<=SIX; digit1<=THREE; digit2<=TWO; digit3<=THREE; end
      16'd3237: begin digit0<=SEVEN; digit1<=THREE; digit2<=TWO; digit3<=THREE; end
      16'd3238: begin digit0<=EIGHT; digit1<=THREE; digit2<=TWO; digit3<=THREE; end
      16'd3239: begin digit0<=NINE; digit1<=THREE; digit2<=TWO; digit3<=THREE; end
      16'd3240: begin digit0<=ZERO; digit1<=FOUR; digit2<=TWO; digit3<=THREE; end
      16'd3241: begin digit0<=ONE; digit1<=FOUR; digit2<=TWO; digit3<=THREE; end
      16'd3242: begin digit0<=TWO; digit1<=FOUR; digit2<=TWO; digit3<=THREE; end
      16'd3243: begin digit0<=THREE; digit1<=FOUR; digit2<=TWO; digit3<=THREE; end
      16'd3244: begin digit0<=FOUR; digit1<=FOUR; digit2<=TWO; digit3<=THREE; end
      16'd3245: begin digit0<=FIVE; digit1<=FOUR; digit2<=TWO; digit3<=THREE; end
      16'd3246: begin digit0<=SIX; digit1<=FOUR; digit2<=TWO; digit3<=THREE; end
      16'd3247: begin digit0<=SEVEN; digit1<=FOUR; digit2<=TWO; digit3<=THREE; end
      16'd3248: begin digit0<=EIGHT; digit1<=FOUR; digit2<=TWO; digit3<=THREE; end
      16'd3249: begin digit0<=NINE; digit1<=FOUR; digit2<=TWO; digit3<=THREE; end
      16'd3250: begin digit0<=ZERO; digit1<=FIVE; digit2<=TWO; digit3<=THREE; end
      16'd3251: begin digit0<=ONE; digit1<=FIVE; digit2<=TWO; digit3<=THREE; end
      16'd3252: begin digit0<=TWO; digit1<=FIVE; digit2<=TWO; digit3<=THREE; end
      16'd3253: begin digit0<=THREE; digit1<=FIVE; digit2<=TWO; digit3<=THREE; end
      16'd3254: begin digit0<=FOUR; digit1<=FIVE; digit2<=TWO; digit3<=THREE; end
      16'd3255: begin digit0<=FIVE; digit1<=FIVE; digit2<=TWO; digit3<=THREE; end
      16'd3256: begin digit0<=SIX; digit1<=FIVE; digit2<=TWO; digit3<=THREE; end
      16'd3257: begin digit0<=SEVEN; digit1<=FIVE; digit2<=TWO; digit3<=THREE; end
      16'd3258: begin digit0<=EIGHT; digit1<=FIVE; digit2<=TWO; digit3<=THREE; end
      16'd3259: begin digit0<=NINE; digit1<=FIVE; digit2<=TWO; digit3<=THREE; end
      16'd3260: begin digit0<=ZERO; digit1<=SIX; digit2<=TWO; digit3<=THREE; end
      16'd3261: begin digit0<=ONE; digit1<=SIX; digit2<=TWO; digit3<=THREE; end
      16'd3262: begin digit0<=TWO; digit1<=SIX; digit2<=TWO; digit3<=THREE; end
      16'd3263: begin digit0<=THREE; digit1<=SIX; digit2<=TWO; digit3<=THREE; end
      16'd3264: begin digit0<=FOUR; digit1<=SIX; digit2<=TWO; digit3<=THREE; end
      16'd3265: begin digit0<=FIVE; digit1<=SIX; digit2<=TWO; digit3<=THREE; end
      16'd3266: begin digit0<=SIX; digit1<=SIX; digit2<=TWO; digit3<=THREE; end
      16'd3267: begin digit0<=SEVEN; digit1<=SIX; digit2<=TWO; digit3<=THREE; end
      16'd3268: begin digit0<=EIGHT; digit1<=SIX; digit2<=TWO; digit3<=THREE; end
      16'd3269: begin digit0<=NINE; digit1<=SIX; digit2<=TWO; digit3<=THREE; end
      16'd3270: begin digit0<=ZERO; digit1<=SEVEN; digit2<=TWO; digit3<=THREE; end
      16'd3271: begin digit0<=ONE; digit1<=SEVEN; digit2<=TWO; digit3<=THREE; end
      16'd3272: begin digit0<=TWO; digit1<=SEVEN; digit2<=TWO; digit3<=THREE; end
      16'd3273: begin digit0<=THREE; digit1<=SEVEN; digit2<=TWO; digit3<=THREE; end
      16'd3274: begin digit0<=FOUR; digit1<=SEVEN; digit2<=TWO; digit3<=THREE; end
      16'd3275: begin digit0<=FIVE; digit1<=SEVEN; digit2<=TWO; digit3<=THREE; end
      16'd3276: begin digit0<=SIX; digit1<=SEVEN; digit2<=TWO; digit3<=THREE; end
      16'd3277: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=TWO; digit3<=THREE; end
      16'd3278: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=TWO; digit3<=THREE; end
      16'd3279: begin digit0<=NINE; digit1<=SEVEN; digit2<=TWO; digit3<=THREE; end
      16'd3280: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=THREE; end
      16'd3281: begin digit0<=ONE; digit1<=EIGHT; digit2<=TWO; digit3<=THREE; end
      16'd3282: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=THREE; end
      16'd3283: begin digit0<=THREE; digit1<=EIGHT; digit2<=TWO; digit3<=THREE; end
      16'd3284: begin digit0<=FOUR; digit1<=EIGHT; digit2<=TWO; digit3<=THREE; end
      16'd3285: begin digit0<=FIVE; digit1<=EIGHT; digit2<=TWO; digit3<=THREE; end
      16'd3286: begin digit0<=SIX; digit1<=EIGHT; digit2<=TWO; digit3<=THREE; end
      16'd3287: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=TWO; digit3<=THREE; end
      16'd3288: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=TWO; digit3<=THREE; end
      16'd3289: begin digit0<=NINE; digit1<=EIGHT; digit2<=TWO; digit3<=THREE; end
      16'd3290: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=THREE; end
      16'd3291: begin digit0<=ONE; digit1<=NINE; digit2<=TWO; digit3<=THREE; end
      16'd3292: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=THREE; end
      16'd3293: begin digit0<=THREE; digit1<=NINE; digit2<=TWO; digit3<=THREE; end
      16'd3294: begin digit0<=FOUR; digit1<=NINE; digit2<=TWO; digit3<=THREE; end
      16'd3295: begin digit0<=FIVE; digit1<=NINE; digit2<=TWO; digit3<=THREE; end
      16'd3296: begin digit0<=SIX; digit1<=NINE; digit2<=TWO; digit3<=THREE; end
      16'd3297: begin digit0<=SEVEN; digit1<=NINE; digit2<=TWO; digit3<=THREE; end
      16'd3298: begin digit0<=EIGHT; digit1<=NINE; digit2<=TWO; digit3<=THREE; end
      16'd3299: begin digit0<=NINE; digit1<=NINE; digit2<=TWO; digit3<=THREE; end
	  16'd3300: begin digit0<=ZERO; digit1<=ZERO; digit2<=THREE; digit3<=THREE; end
      16'd3301: begin digit0<=ONE; digit1<=ZERO; digit2<=THREE; digit3<=THREE; end
      16'd3302: begin digit0<=TWO; digit1<=ZERO; digit2<=THREE; digit3<=THREE; end
      16'd3303: begin digit0<=THREE; digit1<=ZERO; digit2<=THREE; digit3<=THREE; end
      16'd3304: begin digit0<=FOUR; digit1<=ZERO; digit2<=THREE; digit3<=THREE; end
      16'd3305: begin digit0<=FIVE; digit1<=ZERO; digit2<=THREE; digit3<=THREE; end
      16'd3306: begin digit0<=SIX; digit1<=ZERO; digit2<=THREE; digit3<=THREE; end
      16'd3307: begin digit0<=SEVEN; digit1<=ZERO; digit2<=THREE; digit3<=THREE; end
      16'd3308: begin digit0<=EIGHT; digit1<=ZERO; digit2<=THREE; digit3<=THREE; end
      16'd3309: begin digit0<=NINE; digit1<=ZERO; digit2<=THREE; digit3<=THREE; end
      16'd3310: begin digit0<=ZERO; digit1<=ONE; digit2<=THREE; digit3<=THREE; end
      16'd3311: begin digit0<=ONE; digit1<=ONE; digit2<=THREE; digit3<=THREE; end
      16'd3312: begin digit0<=TWO; digit1<=ONE; digit2<=THREE; digit3<=THREE; end
      16'd3313: begin digit0<=THREE; digit1<=ONE; digit2<=THREE; digit3<=THREE; end
      16'd3314: begin digit0<=FOUR; digit1<=ONE; digit2<=THREE; digit3<=THREE; end
      16'd3315: begin digit0<=FIVE; digit1<=ONE; digit2<=THREE; digit3<=THREE; end
      16'd3316: begin digit0<=SIX; digit1<=ONE; digit2<=THREE; digit3<=THREE; end
      16'd3317: begin digit0<=SEVEN; digit1<=ONE; digit2<=THREE; digit3<=THREE; end
      16'd3318: begin digit0<=EIGHT; digit1<=ONE; digit2<=THREE; digit3<=THREE; end
      16'd3319: begin digit0<=NINE; digit1<=ONE; digit2<=THREE; digit3<=THREE; end
      16'd3320: begin digit0<=ZERO; digit1<=TWO; digit2<=THREE; digit3<=THREE; end
      16'd3321: begin digit0<=ONE; digit1<=TWO; digit2<=THREE; digit3<=THREE; end
      16'd3322: begin digit0<=TWO; digit1<=TWO; digit2<=THREE; digit3<=THREE; end
      16'd3323: begin digit0<=THREE; digit1<=TWO; digit2<=THREE; digit3<=THREE; end
      16'd3324: begin digit0<=FOUR; digit1<=TWO; digit2<=THREE; digit3<=THREE; end
      16'd3325: begin digit0<=FIVE; digit1<=TWO; digit2<=THREE; digit3<=THREE; end
      16'd3326: begin digit0<=SIX; digit1<=TWO; digit2<=THREE; digit3<=THREE; end
      16'd3327: begin digit0<=SEVEN; digit1<=TWO; digit2<=THREE; digit3<=THREE; end
      16'd3328: begin digit0<=EIGHT; digit1<=TWO; digit2<=THREE; digit3<=THREE; end
      16'd3329: begin digit0<=NINE; digit1<=TWO; digit2<=THREE; digit3<=THREE; end
      16'd3330: begin digit0<=ZERO; digit1<=THREE; digit2<=THREE; digit3<=THREE; end
      16'd3331: begin digit0<=ONE; digit1<=THREE; digit2<=THREE; digit3<=THREE; end
      16'd3332: begin digit0<=TWO; digit1<=THREE; digit2<=THREE; digit3<=THREE; end
      16'd3333: begin digit0<=THREE; digit1<=THREE; digit2<=THREE; digit3<=THREE; end
      16'd3334: begin digit0<=FOUR; digit1<=THREE; digit2<=THREE; digit3<=THREE; end
      16'd3335: begin digit0<=FIVE; digit1<=THREE; digit2<=THREE; digit3<=THREE; end
      16'd3336: begin digit0<=SIX; digit1<=THREE; digit2<=THREE; digit3<=THREE; end
      16'd3337: begin digit0<=SEVEN; digit1<=THREE; digit2<=THREE; digit3<=THREE; end
      16'd3338: begin digit0<=EIGHT; digit1<=THREE; digit2<=THREE; digit3<=THREE; end
      16'd3339: begin digit0<=NINE; digit1<=THREE; digit2<=THREE; digit3<=THREE; end
      16'd3340: begin digit0<=ZERO; digit1<=FOUR; digit2<=THREE; digit3<=THREE; end
      16'd3341: begin digit0<=ONE; digit1<=FOUR; digit2<=THREE; digit3<=THREE; end
      16'd3342: begin digit0<=TWO; digit1<=FOUR; digit2<=THREE; digit3<=THREE; end
      16'd3343: begin digit0<=THREE; digit1<=FOUR; digit2<=THREE; digit3<=THREE; end
      16'd3344: begin digit0<=FOUR; digit1<=FOUR; digit2<=THREE; digit3<=THREE; end
      16'd3345: begin digit0<=FIVE; digit1<=FOUR; digit2<=THREE; digit3<=THREE; end
      16'd3346: begin digit0<=SIX; digit1<=FOUR; digit2<=THREE; digit3<=THREE; end
      16'd3347: begin digit0<=SEVEN; digit1<=FOUR; digit2<=THREE; digit3<=THREE; end
      16'd3348: begin digit0<=EIGHT; digit1<=FOUR; digit2<=THREE; digit3<=THREE; end
      16'd3349: begin digit0<=NINE; digit1<=FOUR; digit2<=THREE; digit3<=THREE; end
      16'd3350: begin digit0<=ZERO; digit1<=FIVE; digit2<=THREE; digit3<=THREE; end
      16'd3351: begin digit0<=ONE; digit1<=FIVE; digit2<=THREE; digit3<=THREE; end
      16'd3352: begin digit0<=TWO; digit1<=FIVE; digit2<=THREE; digit3<=THREE; end
      16'd3353: begin digit0<=THREE; digit1<=FIVE; digit2<=THREE; digit3<=THREE; end
      16'd3354: begin digit0<=FOUR; digit1<=FIVE; digit2<=THREE; digit3<=THREE; end
      16'd3355: begin digit0<=FIVE; digit1<=FIVE; digit2<=THREE; digit3<=THREE; end
      16'd3356: begin digit0<=SIX; digit1<=FIVE; digit2<=THREE; digit3<=THREE; end
      16'd3357: begin digit0<=SEVEN; digit1<=FIVE; digit2<=THREE; digit3<=THREE; end
      16'd3358: begin digit0<=EIGHT; digit1<=FIVE; digit2<=THREE; digit3<=THREE; end
      16'd3359: begin digit0<=NINE; digit1<=FIVE; digit2<=THREE; digit3<=THREE; end
      16'd3360: begin digit0<=ZERO; digit1<=SIX; digit2<=THREE; digit3<=THREE; end
      16'd3361: begin digit0<=ONE; digit1<=SIX; digit2<=THREE; digit3<=THREE; end
      16'd3362: begin digit0<=TWO; digit1<=SIX; digit2<=THREE; digit3<=THREE; end
      16'd3363: begin digit0<=THREE; digit1<=SIX; digit2<=THREE; digit3<=THREE; end
      16'd3364: begin digit0<=FOUR; digit1<=SIX; digit2<=THREE; digit3<=THREE; end
      16'd3365: begin digit0<=FIVE; digit1<=SIX; digit2<=THREE; digit3<=THREE; end
      16'd3366: begin digit0<=SIX; digit1<=SIX; digit2<=THREE; digit3<=THREE; end
      16'd3367: begin digit0<=SEVEN; digit1<=SIX; digit2<=THREE; digit3<=THREE; end
      16'd3368: begin digit0<=EIGHT; digit1<=SIX; digit2<=THREE; digit3<=THREE; end
      16'd3369: begin digit0<=NINE; digit1<=SIX; digit2<=THREE; digit3<=THREE; end
      16'd3370: begin digit0<=ZERO; digit1<=SEVEN; digit2<=THREE; digit3<=THREE; end
      16'd3371: begin digit0<=ONE; digit1<=SEVEN; digit2<=THREE; digit3<=THREE; end
      16'd3372: begin digit0<=TWO; digit1<=SEVEN; digit2<=THREE; digit3<=THREE; end
      16'd3373: begin digit0<=THREE; digit1<=SEVEN; digit2<=THREE; digit3<=THREE; end
      16'd3374: begin digit0<=FOUR; digit1<=SEVEN; digit2<=THREE; digit3<=THREE; end
      16'd3375: begin digit0<=FIVE; digit1<=SEVEN; digit2<=THREE; digit3<=THREE; end
      16'd3376: begin digit0<=SIX; digit1<=SEVEN; digit2<=THREE; digit3<=THREE; end
      16'd3377: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=THREE; digit3<=THREE; end
      16'd3378: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=THREE; digit3<=THREE; end
      16'd3379: begin digit0<=NINE; digit1<=SEVEN; digit2<=THREE; digit3<=THREE; end
      16'd3380: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=THREE; end
      16'd3381: begin digit0<=ONE; digit1<=EIGHT; digit2<=THREE; digit3<=THREE; end
      16'd3382: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=THREE; end
      16'd3383: begin digit0<=THREE; digit1<=EIGHT; digit2<=THREE; digit3<=THREE; end
      16'd3384: begin digit0<=FOUR; digit1<=EIGHT; digit2<=THREE; digit3<=THREE; end
      16'd3385: begin digit0<=FIVE; digit1<=EIGHT; digit2<=THREE; digit3<=THREE; end
      16'd3386: begin digit0<=SIX; digit1<=EIGHT; digit2<=THREE; digit3<=THREE; end
      16'd3387: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=THREE; digit3<=THREE; end
      16'd3388: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=THREE; digit3<=THREE; end
      16'd3389: begin digit0<=NINE; digit1<=EIGHT; digit2<=THREE; digit3<=THREE; end
      16'd3390: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=THREE; end
      16'd3391: begin digit0<=ONE; digit1<=NINE; digit2<=THREE; digit3<=THREE; end
      16'd3392: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=THREE; end
      16'd3393: begin digit0<=THREE; digit1<=NINE; digit2<=THREE; digit3<=THREE; end
      16'd3394: begin digit0<=FOUR; digit1<=NINE; digit2<=THREE; digit3<=THREE; end
      16'd3395: begin digit0<=FIVE; digit1<=NINE; digit2<=THREE; digit3<=THREE; end
      16'd3396: begin digit0<=SIX; digit1<=NINE; digit2<=THREE; digit3<=THREE; end
      16'd3397: begin digit0<=SEVEN; digit1<=NINE; digit2<=THREE; digit3<=THREE; end
      16'd3398: begin digit0<=EIGHT; digit1<=NINE; digit2<=THREE; digit3<=THREE; end
      16'd3399: begin digit0<=NINE; digit1<=NINE; digit2<=THREE; digit3<=THREE; end
	  16'd3400: begin digit0<=ZERO; digit1<=ZERO; digit2<=FOUR; digit3<=THREE; end
      16'd3401: begin digit0<=ONE; digit1<=ZERO; digit2<=FOUR; digit3<=THREE; end
      16'd3402: begin digit0<=TWO; digit1<=ZERO; digit2<=FOUR; digit3<=THREE; end
      16'd3403: begin digit0<=THREE; digit1<=ZERO; digit2<=FOUR; digit3<=THREE; end
      16'd3404: begin digit0<=FOUR; digit1<=ZERO; digit2<=FOUR; digit3<=THREE; end
      16'd3405: begin digit0<=FIVE; digit1<=ZERO; digit2<=FOUR; digit3<=THREE; end
      16'd3406: begin digit0<=SIX; digit1<=ZERO; digit2<=FOUR; digit3<=THREE; end
      16'd3407: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FOUR; digit3<=THREE; end
      16'd3408: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FOUR; digit3<=THREE; end
      16'd3409: begin digit0<=NINE; digit1<=ZERO; digit2<=FOUR; digit3<=THREE; end
      16'd3410: begin digit0<=ZERO; digit1<=ONE; digit2<=FOUR; digit3<=THREE; end
      16'd3411: begin digit0<=ONE; digit1<=ONE; digit2<=FOUR; digit3<=THREE; end
      16'd3412: begin digit0<=TWO; digit1<=ONE; digit2<=FOUR; digit3<=THREE; end
      16'd3413: begin digit0<=THREE; digit1<=ONE; digit2<=FOUR; digit3<=THREE; end
      16'd3414: begin digit0<=FOUR; digit1<=ONE; digit2<=FOUR; digit3<=THREE; end
      16'd3415: begin digit0<=FIVE; digit1<=ONE; digit2<=FOUR; digit3<=THREE; end
      16'd3416: begin digit0<=SIX; digit1<=ONE; digit2<=FOUR; digit3<=THREE; end
      16'd3417: begin digit0<=SEVEN; digit1<=ONE; digit2<=FOUR; digit3<=THREE; end
      16'd3418: begin digit0<=EIGHT; digit1<=ONE; digit2<=FOUR; digit3<=THREE; end
      16'd3419: begin digit0<=NINE; digit1<=ONE; digit2<=FOUR; digit3<=THREE; end
      16'd3420: begin digit0<=ZERO; digit1<=TWO; digit2<=FOUR; digit3<=THREE; end
      16'd3421: begin digit0<=ONE; digit1<=TWO; digit2<=FOUR; digit3<=THREE; end
      16'd3422: begin digit0<=TWO; digit1<=TWO; digit2<=FOUR; digit3<=THREE; end
      16'd3423: begin digit0<=THREE; digit1<=TWO; digit2<=FOUR; digit3<=THREE; end
      16'd3424: begin digit0<=FOUR; digit1<=TWO; digit2<=FOUR; digit3<=THREE; end
      16'd3425: begin digit0<=FIVE; digit1<=TWO; digit2<=FOUR; digit3<=THREE; end
      16'd3426: begin digit0<=SIX; digit1<=TWO; digit2<=FOUR; digit3<=THREE; end
      16'd3427: begin digit0<=SEVEN; digit1<=TWO; digit2<=FOUR; digit3<=THREE; end
      16'd3428: begin digit0<=EIGHT; digit1<=TWO; digit2<=FOUR; digit3<=THREE; end
      16'd3429: begin digit0<=NINE; digit1<=TWO; digit2<=FOUR; digit3<=THREE; end
      16'd3430: begin digit0<=ZERO; digit1<=THREE; digit2<=FOUR; digit3<=THREE; end
      16'd3431: begin digit0<=ONE; digit1<=THREE; digit2<=FOUR; digit3<=THREE; end
      16'd3432: begin digit0<=TWO; digit1<=THREE; digit2<=FOUR; digit3<=THREE; end
      16'd3433: begin digit0<=THREE; digit1<=THREE; digit2<=FOUR; digit3<=THREE; end
      16'd3434: begin digit0<=FOUR; digit1<=THREE; digit2<=FOUR; digit3<=THREE; end
      16'd3435: begin digit0<=FIVE; digit1<=THREE; digit2<=FOUR; digit3<=THREE; end
      16'd3436: begin digit0<=SIX; digit1<=THREE; digit2<=FOUR; digit3<=THREE; end
      16'd3437: begin digit0<=SEVEN; digit1<=THREE; digit2<=FOUR; digit3<=THREE; end
      16'd3438: begin digit0<=EIGHT; digit1<=THREE; digit2<=FOUR; digit3<=THREE; end
      16'd3439: begin digit0<=NINE; digit1<=THREE; digit2<=FOUR; digit3<=THREE; end
      16'd3440: begin digit0<=ZERO; digit1<=FOUR; digit2<=FOUR; digit3<=THREE; end
      16'd3441: begin digit0<=ONE; digit1<=FOUR; digit2<=FOUR; digit3<=THREE; end
      16'd3442: begin digit0<=TWO; digit1<=FOUR; digit2<=FOUR; digit3<=THREE; end
      16'd3443: begin digit0<=THREE; digit1<=FOUR; digit2<=FOUR; digit3<=THREE; end
      16'd3444: begin digit0<=FOUR; digit1<=FOUR; digit2<=FOUR; digit3<=THREE; end
      16'd3445: begin digit0<=FIVE; digit1<=FOUR; digit2<=FOUR; digit3<=THREE; end
      16'd3446: begin digit0<=SIX; digit1<=FOUR; digit2<=FOUR; digit3<=THREE; end
      16'd3447: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FOUR; digit3<=THREE; end
      16'd3448: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FOUR; digit3<=THREE; end
      16'd3449: begin digit0<=NINE; digit1<=FOUR; digit2<=FOUR; digit3<=THREE; end
      16'd3450: begin digit0<=ZERO; digit1<=FIVE; digit2<=FOUR; digit3<=THREE; end
      16'd3451: begin digit0<=ONE; digit1<=FIVE; digit2<=FOUR; digit3<=THREE; end
      16'd3452: begin digit0<=TWO; digit1<=FIVE; digit2<=FOUR; digit3<=THREE; end
      16'd3453: begin digit0<=THREE; digit1<=FIVE; digit2<=FOUR; digit3<=THREE; end
      16'd3454: begin digit0<=FOUR; digit1<=FIVE; digit2<=FOUR; digit3<=THREE; end
      16'd3455: begin digit0<=FIVE; digit1<=FIVE; digit2<=FOUR; digit3<=THREE; end
      16'd3456: begin digit0<=SIX; digit1<=FIVE; digit2<=FOUR; digit3<=THREE; end
      16'd3457: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FOUR; digit3<=THREE; end
      16'd3458: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FOUR; digit3<=THREE; end
      16'd3459: begin digit0<=NINE; digit1<=FIVE; digit2<=FOUR; digit3<=THREE; end
      16'd3460: begin digit0<=ZERO; digit1<=SIX; digit2<=FOUR; digit3<=THREE; end
      16'd3461: begin digit0<=ONE; digit1<=SIX; digit2<=FOUR; digit3<=THREE; end
      16'd3462: begin digit0<=TWO; digit1<=SIX; digit2<=FOUR; digit3<=THREE; end
      16'd3463: begin digit0<=THREE; digit1<=SIX; digit2<=FOUR; digit3<=THREE; end
      16'd3464: begin digit0<=FOUR; digit1<=SIX; digit2<=FOUR; digit3<=THREE; end
      16'd3465: begin digit0<=FIVE; digit1<=SIX; digit2<=FOUR; digit3<=THREE; end
      16'd3466: begin digit0<=SIX; digit1<=SIX; digit2<=FOUR; digit3<=THREE; end
      16'd3467: begin digit0<=SEVEN; digit1<=SIX; digit2<=FOUR; digit3<=THREE; end
      16'd3468: begin digit0<=EIGHT; digit1<=SIX; digit2<=FOUR; digit3<=THREE; end
      16'd3469: begin digit0<=NINE; digit1<=SIX; digit2<=FOUR; digit3<=THREE; end
      16'd3470: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FOUR; digit3<=THREE; end
      16'd3471: begin digit0<=ONE; digit1<=SEVEN; digit2<=FOUR; digit3<=THREE; end
      16'd3472: begin digit0<=TWO; digit1<=SEVEN; digit2<=FOUR; digit3<=THREE; end
      16'd3473: begin digit0<=THREE; digit1<=SEVEN; digit2<=FOUR; digit3<=THREE; end
      16'd3474: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FOUR; digit3<=THREE; end
      16'd3475: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FOUR; digit3<=THREE; end
      16'd3476: begin digit0<=SIX; digit1<=SEVEN; digit2<=FOUR; digit3<=THREE; end
      16'd3477: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FOUR; digit3<=THREE; end
      16'd3478: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FOUR; digit3<=THREE; end
      16'd3479: begin digit0<=NINE; digit1<=SEVEN; digit2<=FOUR; digit3<=THREE; end
      16'd3480: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=THREE; end
      16'd3481: begin digit0<=ONE; digit1<=EIGHT; digit2<=FOUR; digit3<=THREE; end
      16'd3482: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=THREE; end
      16'd3483: begin digit0<=THREE; digit1<=EIGHT; digit2<=FOUR; digit3<=THREE; end
      16'd3484: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FOUR; digit3<=THREE; end
      16'd3485: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FOUR; digit3<=THREE; end
      16'd3486: begin digit0<=SIX; digit1<=EIGHT; digit2<=FOUR; digit3<=THREE; end
      16'd3487: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FOUR; digit3<=THREE; end
      16'd3488: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FOUR; digit3<=THREE; end
      16'd3489: begin digit0<=NINE; digit1<=EIGHT; digit2<=FOUR; digit3<=THREE; end
      16'd3490: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=THREE; end
      16'd3491: begin digit0<=ONE; digit1<=NINE; digit2<=FOUR; digit3<=THREE; end
      16'd3492: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=THREE; end
      16'd3493: begin digit0<=THREE; digit1<=NINE; digit2<=FOUR; digit3<=THREE; end
      16'd3494: begin digit0<=FOUR; digit1<=NINE; digit2<=FOUR; digit3<=THREE; end
      16'd3495: begin digit0<=FIVE; digit1<=NINE; digit2<=FOUR; digit3<=THREE; end
      16'd3496: begin digit0<=SIX; digit1<=NINE; digit2<=FOUR; digit3<=THREE; end
      16'd3497: begin digit0<=SEVEN; digit1<=NINE; digit2<=FOUR; digit3<=THREE; end
      16'd3498: begin digit0<=EIGHT; digit1<=NINE; digit2<=FOUR; digit3<=THREE; end
      16'd3499: begin digit0<=NINE; digit1<=NINE; digit2<=FOUR; digit3<=THREE; end
	  16'd3500: begin digit0<=ZERO; digit1<=ZERO; digit2<=FIVE; digit3<=THREE; end
      16'd3501: begin digit0<=ONE; digit1<=ZERO; digit2<=FIVE; digit3<=THREE; end
      16'd3502: begin digit0<=TWO; digit1<=ZERO; digit2<=FIVE; digit3<=THREE; end
      16'd3503: begin digit0<=THREE; digit1<=ZERO; digit2<=FIVE; digit3<=THREE; end
      16'd3504: begin digit0<=FOUR; digit1<=ZERO; digit2<=FIVE; digit3<=THREE; end
      16'd3505: begin digit0<=FIVE; digit1<=ZERO; digit2<=FIVE; digit3<=THREE; end
      16'd3506: begin digit0<=SIX; digit1<=ZERO; digit2<=FIVE; digit3<=THREE; end
      16'd3507: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FIVE; digit3<=THREE; end
      16'd3508: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FIVE; digit3<=THREE; end
      16'd3509: begin digit0<=NINE; digit1<=ZERO; digit2<=FIVE; digit3<=THREE; end
      16'd3510: begin digit0<=ZERO; digit1<=ONE; digit2<=FIVE; digit3<=THREE; end
      16'd3511: begin digit0<=ONE; digit1<=ONE; digit2<=FIVE; digit3<=THREE; end
      16'd3512: begin digit0<=TWO; digit1<=ONE; digit2<=FIVE; digit3<=THREE; end
      16'd3513: begin digit0<=THREE; digit1<=ONE; digit2<=FIVE; digit3<=THREE; end
      16'd3514: begin digit0<=FOUR; digit1<=ONE; digit2<=FIVE; digit3<=THREE; end
      16'd3515: begin digit0<=FIVE; digit1<=ONE; digit2<=FIVE; digit3<=THREE; end
      16'd3516: begin digit0<=SIX; digit1<=ONE; digit2<=FIVE; digit3<=THREE; end
      16'd3517: begin digit0<=SEVEN; digit1<=ONE; digit2<=FIVE; digit3<=THREE; end
      16'd3518: begin digit0<=EIGHT; digit1<=ONE; digit2<=FIVE; digit3<=THREE; end
      16'd3519: begin digit0<=NINE; digit1<=ONE; digit2<=FIVE; digit3<=THREE; end
      16'd3520: begin digit0<=ZERO; digit1<=TWO; digit2<=FIVE; digit3<=THREE; end
      16'd3521: begin digit0<=ONE; digit1<=TWO; digit2<=FIVE; digit3<=THREE; end
      16'd3522: begin digit0<=TWO; digit1<=TWO; digit2<=FIVE; digit3<=THREE; end
      16'd3523: begin digit0<=THREE; digit1<=TWO; digit2<=FIVE; digit3<=THREE; end
      16'd3524: begin digit0<=FOUR; digit1<=TWO; digit2<=FIVE; digit3<=THREE; end
      16'd3525: begin digit0<=FIVE; digit1<=TWO; digit2<=FIVE; digit3<=THREE; end
      16'd3526: begin digit0<=SIX; digit1<=TWO; digit2<=FIVE; digit3<=THREE; end
      16'd3527: begin digit0<=SEVEN; digit1<=TWO; digit2<=FIVE; digit3<=THREE; end
      16'd3528: begin digit0<=EIGHT; digit1<=TWO; digit2<=FIVE; digit3<=THREE; end
      16'd3529: begin digit0<=NINE; digit1<=TWO; digit2<=FIVE; digit3<=THREE; end
      16'd3530: begin digit0<=ZERO; digit1<=THREE; digit2<=FIVE; digit3<=THREE; end
      16'd3531: begin digit0<=ONE; digit1<=THREE; digit2<=FIVE; digit3<=THREE; end
      16'd3532: begin digit0<=TWO; digit1<=THREE; digit2<=FIVE; digit3<=THREE; end
      16'd3533: begin digit0<=THREE; digit1<=THREE; digit2<=FIVE; digit3<=THREE; end
      16'd3534: begin digit0<=FOUR; digit1<=THREE; digit2<=FIVE; digit3<=THREE; end
      16'd3535: begin digit0<=FIVE; digit1<=THREE; digit2<=FIVE; digit3<=THREE; end
      16'd3536: begin digit0<=SIX; digit1<=THREE; digit2<=FIVE; digit3<=THREE; end
      16'd3537: begin digit0<=SEVEN; digit1<=THREE; digit2<=FIVE; digit3<=THREE; end
      16'd3538: begin digit0<=EIGHT; digit1<=THREE; digit2<=FIVE; digit3<=THREE; end
      16'd3539: begin digit0<=NINE; digit1<=THREE; digit2<=FIVE; digit3<=THREE; end
      16'd3540: begin digit0<=ZERO; digit1<=FOUR; digit2<=FIVE; digit3<=THREE; end
      16'd3541: begin digit0<=ONE; digit1<=FOUR; digit2<=FIVE; digit3<=THREE; end
      16'd3542: begin digit0<=TWO; digit1<=FOUR; digit2<=FIVE; digit3<=THREE; end
      16'd3543: begin digit0<=THREE; digit1<=FOUR; digit2<=FIVE; digit3<=THREE; end
      16'd3544: begin digit0<=FOUR; digit1<=FOUR; digit2<=FIVE; digit3<=THREE; end
      16'd3545: begin digit0<=FIVE; digit1<=FOUR; digit2<=FIVE; digit3<=THREE; end
      16'd3546: begin digit0<=SIX; digit1<=FOUR; digit2<=FIVE; digit3<=THREE; end
      16'd3547: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FIVE; digit3<=THREE; end
      16'd3548: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FIVE; digit3<=THREE; end
      16'd3549: begin digit0<=NINE; digit1<=FOUR; digit2<=FIVE; digit3<=THREE; end
      16'd3550: begin digit0<=ZERO; digit1<=FIVE; digit2<=FIVE; digit3<=THREE; end
      16'd3551: begin digit0<=ONE; digit1<=FIVE; digit2<=FIVE; digit3<=THREE; end
      16'd3552: begin digit0<=TWO; digit1<=FIVE; digit2<=FIVE; digit3<=THREE; end
      16'd3553: begin digit0<=THREE; digit1<=FIVE; digit2<=FIVE; digit3<=THREE; end
      16'd3554: begin digit0<=FOUR; digit1<=FIVE; digit2<=FIVE; digit3<=THREE; end
      16'd3555: begin digit0<=FIVE; digit1<=FIVE; digit2<=FIVE; digit3<=THREE; end
      16'd3556: begin digit0<=SIX; digit1<=FIVE; digit2<=FIVE; digit3<=THREE; end
      16'd3557: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FIVE; digit3<=THREE; end
      16'd3558: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FIVE; digit3<=THREE; end
      16'd3559: begin digit0<=NINE; digit1<=FIVE; digit2<=FIVE; digit3<=THREE; end
      16'd3560: begin digit0<=ZERO; digit1<=SIX; digit2<=FIVE; digit3<=THREE; end
      16'd3561: begin digit0<=ONE; digit1<=SIX; digit2<=FIVE; digit3<=THREE; end
      16'd3562: begin digit0<=TWO; digit1<=SIX; digit2<=FIVE; digit3<=THREE; end
      16'd3563: begin digit0<=THREE; digit1<=SIX; digit2<=FIVE; digit3<=THREE; end
      16'd3564: begin digit0<=FOUR; digit1<=SIX; digit2<=FIVE; digit3<=THREE; end
      16'd3565: begin digit0<=FIVE; digit1<=SIX; digit2<=FIVE; digit3<=THREE; end
      16'd3566: begin digit0<=SIX; digit1<=SIX; digit2<=FIVE; digit3<=THREE; end
      16'd3567: begin digit0<=SEVEN; digit1<=SIX; digit2<=FIVE; digit3<=THREE; end
      16'd3568: begin digit0<=EIGHT; digit1<=SIX; digit2<=FIVE; digit3<=THREE; end
      16'd3569: begin digit0<=NINE; digit1<=SIX; digit2<=FIVE; digit3<=THREE; end
      16'd3570: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FIVE; digit3<=THREE; end
      16'd3571: begin digit0<=ONE; digit1<=SEVEN; digit2<=FIVE; digit3<=THREE; end
      16'd3572: begin digit0<=TWO; digit1<=SEVEN; digit2<=FIVE; digit3<=THREE; end
      16'd3573: begin digit0<=THREE; digit1<=SEVEN; digit2<=FIVE; digit3<=THREE; end
      16'd3574: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FIVE; digit3<=THREE; end
      16'd3575: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FIVE; digit3<=THREE; end
      16'd3576: begin digit0<=SIX; digit1<=SEVEN; digit2<=FIVE; digit3<=THREE; end
      16'd3577: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FIVE; digit3<=THREE; end
      16'd3578: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FIVE; digit3<=THREE; end
      16'd3579: begin digit0<=NINE; digit1<=SEVEN; digit2<=FIVE; digit3<=THREE; end
      16'd3580: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=THREE; end
      16'd3581: begin digit0<=ONE; digit1<=EIGHT; digit2<=FIVE; digit3<=THREE; end
      16'd3582: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=THREE; end
      16'd3583: begin digit0<=THREE; digit1<=EIGHT; digit2<=FIVE; digit3<=THREE; end
      16'd3584: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FIVE; digit3<=THREE; end
      16'd3585: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FIVE; digit3<=THREE; end
      16'd3586: begin digit0<=SIX; digit1<=EIGHT; digit2<=FIVE; digit3<=THREE; end
      16'd3587: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FIVE; digit3<=THREE; end
      16'd3588: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FIVE; digit3<=THREE; end
      16'd3589: begin digit0<=NINE; digit1<=EIGHT; digit2<=FIVE; digit3<=THREE; end
      16'd3590: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=THREE; end
      16'd3591: begin digit0<=ONE; digit1<=NINE; digit2<=FIVE; digit3<=THREE; end
      16'd3592: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=THREE; end
      16'd3593: begin digit0<=THREE; digit1<=NINE; digit2<=FIVE; digit3<=THREE; end
      16'd3594: begin digit0<=FOUR; digit1<=NINE; digit2<=FIVE; digit3<=THREE; end
      16'd3595: begin digit0<=FIVE; digit1<=NINE; digit2<=FIVE; digit3<=THREE; end
      16'd3596: begin digit0<=SIX; digit1<=NINE; digit2<=FIVE; digit3<=THREE; end
      16'd3597: begin digit0<=SEVEN; digit1<=NINE; digit2<=FIVE; digit3<=THREE; end
      16'd3598: begin digit0<=EIGHT; digit1<=NINE; digit2<=FIVE; digit3<=THREE; end
      16'd3599: begin digit0<=NINE; digit1<=NINE; digit2<=FIVE; digit3<=THREE; end
	  16'd3600: begin digit0<=ZERO; digit1<=ZERO; digit2<=SIX; digit3<=THREE; end
      16'd3601: begin digit0<=ONE; digit1<=ZERO; digit2<=SIX; digit3<=THREE; end
      16'd3602: begin digit0<=TWO; digit1<=ZERO; digit2<=SIX; digit3<=THREE; end
      16'd3603: begin digit0<=THREE; digit1<=ZERO; digit2<=SIX; digit3<=THREE; end
      16'd3604: begin digit0<=FOUR; digit1<=ZERO; digit2<=SIX; digit3<=THREE; end
      16'd3605: begin digit0<=FIVE; digit1<=ZERO; digit2<=SIX; digit3<=THREE; end
      16'd3606: begin digit0<=SIX; digit1<=ZERO; digit2<=SIX; digit3<=THREE; end
      16'd3607: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SIX; digit3<=THREE; end
      16'd3608: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SIX; digit3<=THREE; end
      16'd3609: begin digit0<=NINE; digit1<=ZERO; digit2<=SIX; digit3<=THREE; end
      16'd3610: begin digit0<=ZERO; digit1<=ONE; digit2<=SIX; digit3<=THREE; end
      16'd3611: begin digit0<=ONE; digit1<=ONE; digit2<=SIX; digit3<=THREE; end
      16'd3612: begin digit0<=TWO; digit1<=ONE; digit2<=SIX; digit3<=THREE; end
      16'd3613: begin digit0<=THREE; digit1<=ONE; digit2<=SIX; digit3<=THREE; end
      16'd3614: begin digit0<=FOUR; digit1<=ONE; digit2<=SIX; digit3<=THREE; end
      16'd3615: begin digit0<=FIVE; digit1<=ONE; digit2<=SIX; digit3<=THREE; end
      16'd3616: begin digit0<=SIX; digit1<=ONE; digit2<=SIX; digit3<=THREE; end
      16'd3617: begin digit0<=SEVEN; digit1<=ONE; digit2<=SIX; digit3<=THREE; end
      16'd3618: begin digit0<=EIGHT; digit1<=ONE; digit2<=SIX; digit3<=THREE; end
      16'd3619: begin digit0<=NINE; digit1<=ONE; digit2<=SIX; digit3<=THREE; end
      16'd3620: begin digit0<=ZERO; digit1<=TWO; digit2<=SIX; digit3<=THREE; end
      16'd3621: begin digit0<=ONE; digit1<=TWO; digit2<=SIX; digit3<=THREE; end
      16'd3622: begin digit0<=TWO; digit1<=TWO; digit2<=SIX; digit3<=THREE; end
      16'd3623: begin digit0<=THREE; digit1<=TWO; digit2<=SIX; digit3<=THREE; end
      16'd3624: begin digit0<=FOUR; digit1<=TWO; digit2<=SIX; digit3<=THREE; end
      16'd3625: begin digit0<=FIVE; digit1<=TWO; digit2<=SIX; digit3<=THREE; end
      16'd3626: begin digit0<=SIX; digit1<=TWO; digit2<=SIX; digit3<=THREE; end
      16'd3627: begin digit0<=SEVEN; digit1<=TWO; digit2<=SIX; digit3<=THREE; end
      16'd3628: begin digit0<=EIGHT; digit1<=TWO; digit2<=SIX; digit3<=THREE; end
      16'd3629: begin digit0<=NINE; digit1<=TWO; digit2<=SIX; digit3<=THREE; end
      16'd3630: begin digit0<=ZERO; digit1<=THREE; digit2<=SIX; digit3<=THREE; end
      16'd3631: begin digit0<=ONE; digit1<=THREE; digit2<=SIX; digit3<=THREE; end
      16'd3632: begin digit0<=TWO; digit1<=THREE; digit2<=SIX; digit3<=THREE; end
      16'd3633: begin digit0<=THREE; digit1<=THREE; digit2<=SIX; digit3<=THREE; end
      16'd3634: begin digit0<=FOUR; digit1<=THREE; digit2<=SIX; digit3<=THREE; end
      16'd3635: begin digit0<=FIVE; digit1<=THREE; digit2<=SIX; digit3<=THREE; end
      16'd3636: begin digit0<=SIX; digit1<=THREE; digit2<=SIX; digit3<=THREE; end
      16'd3637: begin digit0<=SEVEN; digit1<=THREE; digit2<=SIX; digit3<=THREE; end
      16'd3638: begin digit0<=EIGHT; digit1<=THREE; digit2<=SIX; digit3<=THREE; end
      16'd3639: begin digit0<=NINE; digit1<=THREE; digit2<=SIX; digit3<=THREE; end
      16'd3640: begin digit0<=ZERO; digit1<=FOUR; digit2<=SIX; digit3<=THREE; end
      16'd3641: begin digit0<=ONE; digit1<=FOUR; digit2<=SIX; digit3<=THREE; end
      16'd3642: begin digit0<=TWO; digit1<=FOUR; digit2<=SIX; digit3<=THREE; end
      16'd3643: begin digit0<=THREE; digit1<=FOUR; digit2<=SIX; digit3<=THREE; end
      16'd3644: begin digit0<=FOUR; digit1<=FOUR; digit2<=SIX; digit3<=THREE; end
      16'd3645: begin digit0<=FIVE; digit1<=FOUR; digit2<=SIX; digit3<=THREE; end
      16'd3646: begin digit0<=SIX; digit1<=FOUR; digit2<=SIX; digit3<=THREE; end
      16'd3647: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SIX; digit3<=THREE; end
      16'd3648: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SIX; digit3<=THREE; end
      16'd3649: begin digit0<=NINE; digit1<=FOUR; digit2<=SIX; digit3<=THREE; end
      16'd3650: begin digit0<=ZERO; digit1<=FIVE; digit2<=SIX; digit3<=THREE; end
      16'd3651: begin digit0<=ONE; digit1<=FIVE; digit2<=SIX; digit3<=THREE; end
      16'd3652: begin digit0<=TWO; digit1<=FIVE; digit2<=SIX; digit3<=THREE; end
      16'd3653: begin digit0<=THREE; digit1<=FIVE; digit2<=SIX; digit3<=THREE; end
      16'd3654: begin digit0<=FOUR; digit1<=FIVE; digit2<=SIX; digit3<=THREE; end
      16'd3655: begin digit0<=FIVE; digit1<=FIVE; digit2<=SIX; digit3<=THREE; end
      16'd3656: begin digit0<=SIX; digit1<=FIVE; digit2<=SIX; digit3<=THREE; end
      16'd3657: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SIX; digit3<=THREE; end
      16'd3658: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SIX; digit3<=THREE; end
      16'd3659: begin digit0<=NINE; digit1<=FIVE; digit2<=SIX; digit3<=THREE; end
      16'd3660: begin digit0<=ZERO; digit1<=SIX; digit2<=SIX; digit3<=THREE; end
      16'd3661: begin digit0<=ONE; digit1<=SIX; digit2<=SIX; digit3<=THREE; end
      16'd3662: begin digit0<=TWO; digit1<=SIX; digit2<=SIX; digit3<=THREE; end
      16'd3663: begin digit0<=THREE; digit1<=SIX; digit2<=SIX; digit3<=THREE; end
      16'd3664: begin digit0<=FOUR; digit1<=SIX; digit2<=SIX; digit3<=THREE; end
      16'd3665: begin digit0<=FIVE; digit1<=SIX; digit2<=SIX; digit3<=THREE; end
      16'd3666: begin digit0<=SIX; digit1<=SIX; digit2<=SIX; digit3<=THREE; end
      16'd3667: begin digit0<=SEVEN; digit1<=SIX; digit2<=SIX; digit3<=THREE; end
      16'd3668: begin digit0<=EIGHT; digit1<=SIX; digit2<=SIX; digit3<=THREE; end
      16'd3669: begin digit0<=NINE; digit1<=SIX; digit2<=SIX; digit3<=THREE; end
      16'd3670: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SIX; digit3<=THREE; end
      16'd3671: begin digit0<=ONE; digit1<=SEVEN; digit2<=SIX; digit3<=THREE; end
      16'd3672: begin digit0<=TWO; digit1<=SEVEN; digit2<=SIX; digit3<=THREE; end
      16'd3673: begin digit0<=THREE; digit1<=SEVEN; digit2<=SIX; digit3<=THREE; end
      16'd3674: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SIX; digit3<=THREE; end
      16'd3675: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SIX; digit3<=THREE; end
      16'd3676: begin digit0<=SIX; digit1<=SEVEN; digit2<=SIX; digit3<=THREE; end
      16'd3677: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SIX; digit3<=THREE; end
      16'd3678: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SIX; digit3<=THREE; end
      16'd3679: begin digit0<=NINE; digit1<=SEVEN; digit2<=SIX; digit3<=THREE; end
      16'd3680: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=THREE; end
      16'd3681: begin digit0<=ONE; digit1<=EIGHT; digit2<=SIX; digit3<=THREE; end
      16'd3682: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=THREE; end
      16'd3683: begin digit0<=THREE; digit1<=EIGHT; digit2<=SIX; digit3<=THREE; end
      16'd3684: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SIX; digit3<=THREE; end
      16'd3685: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SIX; digit3<=THREE; end
      16'd3686: begin digit0<=SIX; digit1<=EIGHT; digit2<=SIX; digit3<=THREE; end
      16'd3687: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SIX; digit3<=THREE; end
      16'd3688: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SIX; digit3<=THREE; end
      16'd3689: begin digit0<=NINE; digit1<=EIGHT; digit2<=SIX; digit3<=THREE; end
      16'd3690: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=THREE; end
      16'd3691: begin digit0<=ONE; digit1<=NINE; digit2<=SIX; digit3<=THREE; end
      16'd3692: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=THREE; end
      16'd3693: begin digit0<=THREE; digit1<=NINE; digit2<=SIX; digit3<=THREE; end
      16'd3694: begin digit0<=FOUR; digit1<=NINE; digit2<=SIX; digit3<=THREE; end
      16'd3695: begin digit0<=FIVE; digit1<=NINE; digit2<=SIX; digit3<=THREE; end
      16'd3696: begin digit0<=SIX; digit1<=NINE; digit2<=SIX; digit3<=THREE; end
      16'd3697: begin digit0<=SEVEN; digit1<=NINE; digit2<=SIX; digit3<=THREE; end
      16'd3698: begin digit0<=EIGHT; digit1<=NINE; digit2<=SIX; digit3<=THREE; end
      16'd3699: begin digit0<=NINE; digit1<=NINE; digit2<=SIX; digit3<=THREE; end
	  16'd3700: begin digit0<=ZERO; digit1<=ZERO; digit2<=SEVEN; digit3<=THREE; end
      16'd3701: begin digit0<=ONE; digit1<=ZERO; digit2<=SEVEN; digit3<=THREE; end
      16'd3702: begin digit0<=TWO; digit1<=ZERO; digit2<=SEVEN; digit3<=THREE; end
      16'd3703: begin digit0<=THREE; digit1<=ZERO; digit2<=SEVEN; digit3<=THREE; end
      16'd3704: begin digit0<=FOUR; digit1<=ZERO; digit2<=SEVEN; digit3<=THREE; end
      16'd3705: begin digit0<=FIVE; digit1<=ZERO; digit2<=SEVEN; digit3<=THREE; end
      16'd3706: begin digit0<=SIX; digit1<=ZERO; digit2<=SEVEN; digit3<=THREE; end
      16'd3707: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SEVEN; digit3<=THREE; end
      16'd3708: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SEVEN; digit3<=THREE; end
      16'd3709: begin digit0<=NINE; digit1<=ZERO; digit2<=SEVEN; digit3<=THREE; end
      16'd3710: begin digit0<=ZERO; digit1<=ONE; digit2<=SEVEN; digit3<=THREE; end
      16'd3711: begin digit0<=ONE; digit1<=ONE; digit2<=SEVEN; digit3<=THREE; end
      16'd3712: begin digit0<=TWO; digit1<=ONE; digit2<=SEVEN; digit3<=THREE; end
      16'd3713: begin digit0<=THREE; digit1<=ONE; digit2<=SEVEN; digit3<=THREE; end
      16'd3714: begin digit0<=FOUR; digit1<=ONE; digit2<=SEVEN; digit3<=THREE; end
      16'd3715: begin digit0<=FIVE; digit1<=ONE; digit2<=SEVEN; digit3<=THREE; end
      16'd3716: begin digit0<=SIX; digit1<=ONE; digit2<=SEVEN; digit3<=THREE; end
      16'd3717: begin digit0<=SEVEN; digit1<=ONE; digit2<=SEVEN; digit3<=THREE; end
      16'd3718: begin digit0<=EIGHT; digit1<=ONE; digit2<=SEVEN; digit3<=THREE; end
      16'd3719: begin digit0<=NINE; digit1<=ONE; digit2<=SEVEN; digit3<=THREE; end
      16'd3720: begin digit0<=ZERO; digit1<=TWO; digit2<=SEVEN; digit3<=THREE; end
      16'd3721: begin digit0<=ONE; digit1<=TWO; digit2<=SEVEN; digit3<=THREE; end
      16'd3722: begin digit0<=TWO; digit1<=TWO; digit2<=SEVEN; digit3<=THREE; end
      16'd3723: begin digit0<=THREE; digit1<=TWO; digit2<=SEVEN; digit3<=THREE; end
      16'd3724: begin digit0<=FOUR; digit1<=TWO; digit2<=SEVEN; digit3<=THREE; end
      16'd3725: begin digit0<=FIVE; digit1<=TWO; digit2<=SEVEN; digit3<=THREE; end
      16'd3726: begin digit0<=SIX; digit1<=TWO; digit2<=SEVEN; digit3<=THREE; end
      16'd3727: begin digit0<=SEVEN; digit1<=TWO; digit2<=SEVEN; digit3<=THREE; end
      16'd3728: begin digit0<=EIGHT; digit1<=TWO; digit2<=SEVEN; digit3<=THREE; end
      16'd3729: begin digit0<=NINE; digit1<=TWO; digit2<=SEVEN; digit3<=THREE; end
      16'd3730: begin digit0<=ZERO; digit1<=THREE; digit2<=SEVEN; digit3<=THREE; end
      16'd3731: begin digit0<=ONE; digit1<=THREE; digit2<=SEVEN; digit3<=THREE; end
      16'd3732: begin digit0<=TWO; digit1<=THREE; digit2<=SEVEN; digit3<=THREE; end
      16'd3733: begin digit0<=THREE; digit1<=THREE; digit2<=SEVEN; digit3<=THREE; end
      16'd3734: begin digit0<=FOUR; digit1<=THREE; digit2<=SEVEN; digit3<=THREE; end
      16'd3735: begin digit0<=FIVE; digit1<=THREE; digit2<=SEVEN; digit3<=THREE; end
      16'd3736: begin digit0<=SIX; digit1<=THREE; digit2<=SEVEN; digit3<=THREE; end
      16'd3737: begin digit0<=SEVEN; digit1<=THREE; digit2<=SEVEN; digit3<=THREE; end
      16'd3738: begin digit0<=EIGHT; digit1<=THREE; digit2<=SEVEN; digit3<=THREE; end
      16'd3739: begin digit0<=NINE; digit1<=THREE; digit2<=SEVEN; digit3<=THREE; end
      16'd3740: begin digit0<=ZERO; digit1<=FOUR; digit2<=SEVEN; digit3<=THREE; end
      16'd3741: begin digit0<=ONE; digit1<=FOUR; digit2<=SEVEN; digit3<=THREE; end
      16'd3742: begin digit0<=TWO; digit1<=FOUR; digit2<=SEVEN; digit3<=THREE; end
      16'd3743: begin digit0<=THREE; digit1<=FOUR; digit2<=SEVEN; digit3<=THREE; end
      16'd3744: begin digit0<=FOUR; digit1<=FOUR; digit2<=SEVEN; digit3<=THREE; end
      16'd3745: begin digit0<=FIVE; digit1<=FOUR; digit2<=SEVEN; digit3<=THREE; end
      16'd3746: begin digit0<=SIX; digit1<=FOUR; digit2<=SEVEN; digit3<=THREE; end
      16'd3747: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SEVEN; digit3<=THREE; end
      16'd3748: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SEVEN; digit3<=THREE; end
      16'd3749: begin digit0<=NINE; digit1<=FOUR; digit2<=SEVEN; digit3<=THREE; end
      16'd3750: begin digit0<=ZERO; digit1<=FIVE; digit2<=SEVEN; digit3<=THREE; end
      16'd3751: begin digit0<=ONE; digit1<=FIVE; digit2<=SEVEN; digit3<=THREE; end
      16'd3752: begin digit0<=TWO; digit1<=FIVE; digit2<=SEVEN; digit3<=THREE; end
      16'd3753: begin digit0<=THREE; digit1<=FIVE; digit2<=SEVEN; digit3<=THREE; end
      16'd3754: begin digit0<=FOUR; digit1<=FIVE; digit2<=SEVEN; digit3<=THREE; end
      16'd3755: begin digit0<=FIVE; digit1<=FIVE; digit2<=SEVEN; digit3<=THREE; end
      16'd3756: begin digit0<=SIX; digit1<=FIVE; digit2<=SEVEN; digit3<=THREE; end
      16'd3757: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SEVEN; digit3<=THREE; end
      16'd3758: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SEVEN; digit3<=THREE; end
      16'd3759: begin digit0<=NINE; digit1<=FIVE; digit2<=SEVEN; digit3<=THREE; end
      16'd3760: begin digit0<=ZERO; digit1<=SIX; digit2<=SEVEN; digit3<=THREE; end
      16'd3761: begin digit0<=ONE; digit1<=SIX; digit2<=SEVEN; digit3<=THREE; end
      16'd3762: begin digit0<=TWO; digit1<=SIX; digit2<=SEVEN; digit3<=THREE; end
      16'd3763: begin digit0<=THREE; digit1<=SIX; digit2<=SEVEN; digit3<=THREE; end
      16'd3764: begin digit0<=FOUR; digit1<=SIX; digit2<=SEVEN; digit3<=THREE; end
      16'd3765: begin digit0<=FIVE; digit1<=SIX; digit2<=SEVEN; digit3<=THREE; end
      16'd3766: begin digit0<=SIX; digit1<=SIX; digit2<=SEVEN; digit3<=THREE; end
      16'd3767: begin digit0<=SEVEN; digit1<=SIX; digit2<=SEVEN; digit3<=THREE; end
      16'd3768: begin digit0<=EIGHT; digit1<=SIX; digit2<=SEVEN; digit3<=THREE; end
      16'd3769: begin digit0<=NINE; digit1<=SIX; digit2<=SEVEN; digit3<=THREE; end
      16'd3770: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SEVEN; digit3<=THREE; end
      16'd3771: begin digit0<=ONE; digit1<=SEVEN; digit2<=SEVEN; digit3<=THREE; end
      16'd3772: begin digit0<=TWO; digit1<=SEVEN; digit2<=SEVEN; digit3<=THREE; end
      16'd3773: begin digit0<=THREE; digit1<=SEVEN; digit2<=SEVEN; digit3<=THREE; end
      16'd3774: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SEVEN; digit3<=THREE; end
      16'd3775: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SEVEN; digit3<=THREE; end
      16'd3776: begin digit0<=SIX; digit1<=SEVEN; digit2<=SEVEN; digit3<=THREE; end
      16'd3777: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SEVEN; digit3<=THREE; end
      16'd3778: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SEVEN; digit3<=THREE; end
      16'd3779: begin digit0<=NINE; digit1<=SEVEN; digit2<=SEVEN; digit3<=THREE; end
      16'd3780: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=THREE; end
      16'd3781: begin digit0<=ONE; digit1<=EIGHT; digit2<=SEVEN; digit3<=THREE; end
      16'd3782: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=THREE; end
      16'd3783: begin digit0<=THREE; digit1<=EIGHT; digit2<=SEVEN; digit3<=THREE; end
      16'd3784: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SEVEN; digit3<=THREE; end
      16'd3785: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SEVEN; digit3<=THREE; end
      16'd3786: begin digit0<=SIX; digit1<=EIGHT; digit2<=SEVEN; digit3<=THREE; end
      16'd3787: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SEVEN; digit3<=THREE; end
      16'd3788: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SEVEN; digit3<=THREE; end
      16'd3789: begin digit0<=NINE; digit1<=EIGHT; digit2<=SEVEN; digit3<=THREE; end
      16'd3790: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=THREE; end
      16'd3791: begin digit0<=ONE; digit1<=NINE; digit2<=SEVEN; digit3<=THREE; end
      16'd3792: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=THREE; end
      16'd3793: begin digit0<=THREE; digit1<=NINE; digit2<=SEVEN; digit3<=THREE; end
      16'd3794: begin digit0<=FOUR; digit1<=NINE; digit2<=SEVEN; digit3<=THREE; end
      16'd3795: begin digit0<=FIVE; digit1<=NINE; digit2<=SEVEN; digit3<=THREE; end
      16'd3796: begin digit0<=SIX; digit1<=NINE; digit2<=SEVEN; digit3<=THREE; end
      16'd3797: begin digit0<=SEVEN; digit1<=NINE; digit2<=SEVEN; digit3<=THREE; end
      16'd3798: begin digit0<=EIGHT; digit1<=NINE; digit2<=SEVEN; digit3<=THREE; end
      16'd3799: begin digit0<=NINE; digit1<=NINE; digit2<=SEVEN; digit3<=THREE; end
	  16'd3800: begin digit0<=ZERO; digit1<=ZERO; digit2<=EIGHT; digit3<=THREE; end
      16'd3801: begin digit0<=ONE; digit1<=ZERO; digit2<=EIGHT; digit3<=THREE; end
      16'd3802: begin digit0<=TWO; digit1<=ZERO; digit2<=EIGHT; digit3<=THREE; end
      16'd3803: begin digit0<=THREE; digit1<=ZERO; digit2<=EIGHT; digit3<=THREE; end
      16'd3804: begin digit0<=FOUR; digit1<=ZERO; digit2<=EIGHT; digit3<=THREE; end
      16'd3805: begin digit0<=FIVE; digit1<=ZERO; digit2<=EIGHT; digit3<=THREE; end
      16'd3806: begin digit0<=SIX; digit1<=ZERO; digit2<=EIGHT; digit3<=THREE; end
      16'd3807: begin digit0<=SEVEN; digit1<=ZERO; digit2<=EIGHT; digit3<=THREE; end
      16'd3808: begin digit0<=EIGHT; digit1<=ZERO; digit2<=EIGHT; digit3<=THREE; end
      16'd3809: begin digit0<=NINE; digit1<=ZERO; digit2<=EIGHT; digit3<=THREE; end
      16'd3810: begin digit0<=ZERO; digit1<=ONE; digit2<=EIGHT; digit3<=THREE; end
      16'd3811: begin digit0<=ONE; digit1<=ONE; digit2<=EIGHT; digit3<=THREE; end
      16'd3812: begin digit0<=TWO; digit1<=ONE; digit2<=EIGHT; digit3<=THREE; end
      16'd3813: begin digit0<=THREE; digit1<=ONE; digit2<=EIGHT; digit3<=THREE; end
      16'd3814: begin digit0<=FOUR; digit1<=ONE; digit2<=EIGHT; digit3<=THREE; end
      16'd3815: begin digit0<=FIVE; digit1<=ONE; digit2<=EIGHT; digit3<=THREE; end
      16'd3816: begin digit0<=SIX; digit1<=ONE; digit2<=EIGHT; digit3<=THREE; end
      16'd3817: begin digit0<=SEVEN; digit1<=ONE; digit2<=EIGHT; digit3<=THREE; end
      16'd3818: begin digit0<=EIGHT; digit1<=ONE; digit2<=EIGHT; digit3<=THREE; end
      16'd3819: begin digit0<=NINE; digit1<=ONE; digit2<=EIGHT; digit3<=THREE; end
      16'd3820: begin digit0<=ZERO; digit1<=TWO; digit2<=EIGHT; digit3<=THREE; end
      16'd3821: begin digit0<=ONE; digit1<=TWO; digit2<=EIGHT; digit3<=THREE; end
      16'd3822: begin digit0<=TWO; digit1<=TWO; digit2<=EIGHT; digit3<=THREE; end
      16'd3823: begin digit0<=THREE; digit1<=TWO; digit2<=EIGHT; digit3<=THREE; end
      16'd3824: begin digit0<=FOUR; digit1<=TWO; digit2<=EIGHT; digit3<=THREE; end
      16'd3825: begin digit0<=FIVE; digit1<=TWO; digit2<=EIGHT; digit3<=THREE; end
      16'd3826: begin digit0<=SIX; digit1<=TWO; digit2<=EIGHT; digit3<=THREE; end
      16'd3827: begin digit0<=SEVEN; digit1<=TWO; digit2<=EIGHT; digit3<=THREE; end
      16'd3828: begin digit0<=EIGHT; digit1<=TWO; digit2<=EIGHT; digit3<=THREE; end
      16'd3829: begin digit0<=NINE; digit1<=TWO; digit2<=EIGHT; digit3<=THREE; end
      16'd3830: begin digit0<=ZERO; digit1<=THREE; digit2<=EIGHT; digit3<=THREE; end
      16'd3831: begin digit0<=ONE; digit1<=THREE; digit2<=EIGHT; digit3<=THREE; end
      16'd3832: begin digit0<=TWO; digit1<=THREE; digit2<=EIGHT; digit3<=THREE; end
      16'd3833: begin digit0<=THREE; digit1<=THREE; digit2<=EIGHT; digit3<=THREE; end
      16'd3834: begin digit0<=FOUR; digit1<=THREE; digit2<=EIGHT; digit3<=THREE; end
      16'd3835: begin digit0<=FIVE; digit1<=THREE; digit2<=EIGHT; digit3<=THREE; end
      16'd3836: begin digit0<=SIX; digit1<=THREE; digit2<=EIGHT; digit3<=THREE; end
      16'd3837: begin digit0<=SEVEN; digit1<=THREE; digit2<=EIGHT; digit3<=THREE; end
      16'd3838: begin digit0<=EIGHT; digit1<=THREE; digit2<=EIGHT; digit3<=THREE; end
      16'd3839: begin digit0<=NINE; digit1<=THREE; digit2<=EIGHT; digit3<=THREE; end
      16'd3840: begin digit0<=ZERO; digit1<=FOUR; digit2<=EIGHT; digit3<=THREE; end
      16'd3841: begin digit0<=ONE; digit1<=FOUR; digit2<=EIGHT; digit3<=THREE; end
      16'd3842: begin digit0<=TWO; digit1<=FOUR; digit2<=EIGHT; digit3<=THREE; end
      16'd3843: begin digit0<=THREE; digit1<=FOUR; digit2<=EIGHT; digit3<=THREE; end
      16'd3844: begin digit0<=FOUR; digit1<=FOUR; digit2<=EIGHT; digit3<=THREE; end
      16'd3845: begin digit0<=FIVE; digit1<=FOUR; digit2<=EIGHT; digit3<=THREE; end
      16'd3846: begin digit0<=SIX; digit1<=FOUR; digit2<=EIGHT; digit3<=THREE; end
      16'd3847: begin digit0<=SEVEN; digit1<=FOUR; digit2<=EIGHT; digit3<=THREE; end
      16'd3848: begin digit0<=EIGHT; digit1<=FOUR; digit2<=EIGHT; digit3<=THREE; end
      16'd3849: begin digit0<=NINE; digit1<=FOUR; digit2<=EIGHT; digit3<=THREE; end
      16'd3850: begin digit0<=ZERO; digit1<=FIVE; digit2<=EIGHT; digit3<=THREE; end
      16'd3851: begin digit0<=ONE; digit1<=FIVE; digit2<=EIGHT; digit3<=THREE; end
      16'd3852: begin digit0<=TWO; digit1<=FIVE; digit2<=EIGHT; digit3<=THREE; end
      16'd3853: begin digit0<=THREE; digit1<=FIVE; digit2<=EIGHT; digit3<=THREE; end
      16'd3854: begin digit0<=FOUR; digit1<=FIVE; digit2<=EIGHT; digit3<=THREE; end
      16'd3855: begin digit0<=FIVE; digit1<=FIVE; digit2<=EIGHT; digit3<=THREE; end
      16'd3856: begin digit0<=SIX; digit1<=FIVE; digit2<=EIGHT; digit3<=THREE; end
      16'd3857: begin digit0<=SEVEN; digit1<=FIVE; digit2<=EIGHT; digit3<=THREE; end
      16'd3858: begin digit0<=EIGHT; digit1<=FIVE; digit2<=EIGHT; digit3<=THREE; end
      16'd3859: begin digit0<=NINE; digit1<=FIVE; digit2<=EIGHT; digit3<=THREE; end
      16'd3860: begin digit0<=ZERO; digit1<=SIX; digit2<=EIGHT; digit3<=THREE; end
      16'd3861: begin digit0<=ONE; digit1<=SIX; digit2<=EIGHT; digit3<=THREE; end
      16'd3862: begin digit0<=TWO; digit1<=SIX; digit2<=EIGHT; digit3<=THREE; end
      16'd3863: begin digit0<=THREE; digit1<=SIX; digit2<=EIGHT; digit3<=THREE; end
      16'd3864: begin digit0<=FOUR; digit1<=SIX; digit2<=EIGHT; digit3<=THREE; end
      16'd3865: begin digit0<=FIVE; digit1<=SIX; digit2<=EIGHT; digit3<=THREE; end
      16'd3866: begin digit0<=SIX; digit1<=SIX; digit2<=EIGHT; digit3<=THREE; end
      16'd3867: begin digit0<=SEVEN; digit1<=SIX; digit2<=EIGHT; digit3<=THREE; end
      16'd3868: begin digit0<=EIGHT; digit1<=SIX; digit2<=EIGHT; digit3<=THREE; end
      16'd3869: begin digit0<=NINE; digit1<=SIX; digit2<=EIGHT; digit3<=THREE; end
      16'd3870: begin digit0<=ZERO; digit1<=SEVEN; digit2<=EIGHT; digit3<=THREE; end
      16'd3871: begin digit0<=ONE; digit1<=SEVEN; digit2<=EIGHT; digit3<=THREE; end
      16'd3872: begin digit0<=TWO; digit1<=SEVEN; digit2<=EIGHT; digit3<=THREE; end
      16'd3873: begin digit0<=THREE; digit1<=SEVEN; digit2<=EIGHT; digit3<=THREE; end
      16'd3874: begin digit0<=FOUR; digit1<=SEVEN; digit2<=EIGHT; digit3<=THREE; end
      16'd3875: begin digit0<=FIVE; digit1<=SEVEN; digit2<=EIGHT; digit3<=THREE; end
      16'd3876: begin digit0<=SIX; digit1<=SEVEN; digit2<=EIGHT; digit3<=THREE; end
      16'd3877: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=EIGHT; digit3<=THREE; end
      16'd3878: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=EIGHT; digit3<=THREE; end
      16'd3879: begin digit0<=NINE; digit1<=SEVEN; digit2<=EIGHT; digit3<=THREE; end
      16'd3880: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=THREE; end
      16'd3881: begin digit0<=ONE; digit1<=EIGHT; digit2<=EIGHT; digit3<=THREE; end
      16'd3882: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=THREE; end
      16'd3883: begin digit0<=THREE; digit1<=EIGHT; digit2<=EIGHT; digit3<=THREE; end
      16'd3884: begin digit0<=FOUR; digit1<=EIGHT; digit2<=EIGHT; digit3<=THREE; end
      16'd3885: begin digit0<=FIVE; digit1<=EIGHT; digit2<=EIGHT; digit3<=THREE; end
      16'd3886: begin digit0<=SIX; digit1<=EIGHT; digit2<=EIGHT; digit3<=THREE; end
      16'd3887: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=EIGHT; digit3<=THREE; end
      16'd3888: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=EIGHT; digit3<=THREE; end
      16'd3889: begin digit0<=NINE; digit1<=EIGHT; digit2<=EIGHT; digit3<=THREE; end
      16'd3890: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=THREE; end
      16'd3891: begin digit0<=ONE; digit1<=NINE; digit2<=EIGHT; digit3<=THREE; end
      16'd3892: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=THREE; end
      16'd3893: begin digit0<=THREE; digit1<=NINE; digit2<=EIGHT; digit3<=THREE; end
      16'd3894: begin digit0<=FOUR; digit1<=NINE; digit2<=EIGHT; digit3<=THREE; end
      16'd3895: begin digit0<=FIVE; digit1<=NINE; digit2<=EIGHT; digit3<=THREE; end
      16'd3896: begin digit0<=SIX; digit1<=NINE; digit2<=EIGHT; digit3<=THREE; end
      16'd3897: begin digit0<=SEVEN; digit1<=NINE; digit2<=EIGHT; digit3<=THREE; end
      16'd3898: begin digit0<=EIGHT; digit1<=NINE; digit2<=EIGHT; digit3<=THREE; end
      16'd3899: begin digit0<=NINE; digit1<=NINE; digit2<=EIGHT; digit3<=THREE; end
	  16'd3900: begin digit0<=ZERO; digit1<=ZERO; digit2<=NINE; digit3<=THREE; end
      16'd3901: begin digit0<=ONE; digit1<=ZERO; digit2<=NINE; digit3<=THREE; end
      16'd3902: begin digit0<=TWO; digit1<=ZERO; digit2<=NINE; digit3<=THREE; end
      16'd3903: begin digit0<=THREE; digit1<=ZERO; digit2<=NINE; digit3<=THREE; end
      16'd3904: begin digit0<=FOUR; digit1<=ZERO; digit2<=NINE; digit3<=THREE; end
      16'd3905: begin digit0<=FIVE; digit1<=ZERO; digit2<=NINE; digit3<=THREE; end
      16'd3906: begin digit0<=SIX; digit1<=ZERO; digit2<=NINE; digit3<=THREE; end
      16'd3907: begin digit0<=SEVEN; digit1<=ZERO; digit2<=NINE; digit3<=THREE; end
      16'd3908: begin digit0<=EIGHT; digit1<=ZERO; digit2<=NINE; digit3<=THREE; end
      16'd3909: begin digit0<=NINE; digit1<=ZERO; digit2<=NINE; digit3<=THREE; end
      16'd3910: begin digit0<=ZERO; digit1<=ONE; digit2<=NINE; digit3<=THREE; end
      16'd3911: begin digit0<=ONE; digit1<=ONE; digit2<=NINE; digit3<=THREE; end
      16'd3912: begin digit0<=TWO; digit1<=ONE; digit2<=NINE; digit3<=THREE; end
      16'd3913: begin digit0<=THREE; digit1<=ONE; digit2<=NINE; digit3<=THREE; end
      16'd3914: begin digit0<=FOUR; digit1<=ONE; digit2<=NINE; digit3<=THREE; end
      16'd3915: begin digit0<=FIVE; digit1<=ONE; digit2<=NINE; digit3<=THREE; end
      16'd3916: begin digit0<=SIX; digit1<=ONE; digit2<=NINE; digit3<=THREE; end
      16'd3917: begin digit0<=SEVEN; digit1<=ONE; digit2<=NINE; digit3<=THREE; end
      16'd3918: begin digit0<=EIGHT; digit1<=ONE; digit2<=NINE; digit3<=THREE; end
      16'd3919: begin digit0<=NINE; digit1<=ONE; digit2<=NINE; digit3<=THREE; end
      16'd3920: begin digit0<=ZERO; digit1<=TWO; digit2<=NINE; digit3<=THREE; end
      16'd3921: begin digit0<=ONE; digit1<=TWO; digit2<=NINE; digit3<=THREE; end
      16'd3922: begin digit0<=TWO; digit1<=TWO; digit2<=NINE; digit3<=THREE; end
      16'd3923: begin digit0<=THREE; digit1<=TWO; digit2<=NINE; digit3<=THREE; end
      16'd3924: begin digit0<=FOUR; digit1<=TWO; digit2<=NINE; digit3<=THREE; end
      16'd3925: begin digit0<=FIVE; digit1<=TWO; digit2<=NINE; digit3<=THREE; end
      16'd3926: begin digit0<=SIX; digit1<=TWO; digit2<=NINE; digit3<=THREE; end
      16'd3927: begin digit0<=SEVEN; digit1<=TWO; digit2<=NINE; digit3<=THREE; end
      16'd3928: begin digit0<=EIGHT; digit1<=TWO; digit2<=NINE; digit3<=THREE; end
      16'd3929: begin digit0<=NINE; digit1<=TWO; digit2<=NINE; digit3<=THREE; end
      16'd3930: begin digit0<=ZERO; digit1<=THREE; digit2<=NINE; digit3<=THREE; end
      16'd3931: begin digit0<=ONE; digit1<=THREE; digit2<=NINE; digit3<=THREE; end
      16'd3932: begin digit0<=TWO; digit1<=THREE; digit2<=NINE; digit3<=THREE; end
      16'd3933: begin digit0<=THREE; digit1<=THREE; digit2<=NINE; digit3<=THREE; end
      16'd3934: begin digit0<=FOUR; digit1<=THREE; digit2<=NINE; digit3<=THREE; end
      16'd3935: begin digit0<=FIVE; digit1<=THREE; digit2<=NINE; digit3<=THREE; end
      16'd3936: begin digit0<=SIX; digit1<=THREE; digit2<=NINE; digit3<=THREE; end
      16'd3937: begin digit0<=SEVEN; digit1<=THREE; digit2<=NINE; digit3<=THREE; end
      16'd3938: begin digit0<=EIGHT; digit1<=THREE; digit2<=NINE; digit3<=THREE; end
      16'd3939: begin digit0<=NINE; digit1<=THREE; digit2<=NINE; digit3<=THREE; end
      16'd3940: begin digit0<=ZERO; digit1<=FOUR; digit2<=NINE; digit3<=THREE; end
      16'd3941: begin digit0<=ONE; digit1<=FOUR; digit2<=NINE; digit3<=THREE; end
      16'd3942: begin digit0<=TWO; digit1<=FOUR; digit2<=NINE; digit3<=THREE; end
      16'd3943: begin digit0<=THREE; digit1<=FOUR; digit2<=NINE; digit3<=THREE; end
      16'd3944: begin digit0<=FOUR; digit1<=FOUR; digit2<=NINE; digit3<=THREE; end
      16'd3945: begin digit0<=FIVE; digit1<=FOUR; digit2<=NINE; digit3<=THREE; end
      16'd3946: begin digit0<=SIX; digit1<=FOUR; digit2<=NINE; digit3<=THREE; end
      16'd3947: begin digit0<=SEVEN; digit1<=FOUR; digit2<=NINE; digit3<=THREE; end
      16'd3948: begin digit0<=EIGHT; digit1<=FOUR; digit2<=NINE; digit3<=THREE; end
      16'd3949: begin digit0<=NINE; digit1<=FOUR; digit2<=NINE; digit3<=THREE; end
      16'd3950: begin digit0<=ZERO; digit1<=FIVE; digit2<=NINE; digit3<=THREE; end
      16'd3951: begin digit0<=ONE; digit1<=FIVE; digit2<=NINE; digit3<=THREE; end
      16'd3952: begin digit0<=TWO; digit1<=FIVE; digit2<=NINE; digit3<=THREE; end
      16'd3953: begin digit0<=THREE; digit1<=FIVE; digit2<=NINE; digit3<=THREE; end
      16'd3954: begin digit0<=FOUR; digit1<=FIVE; digit2<=NINE; digit3<=THREE; end
      16'd3955: begin digit0<=FIVE; digit1<=FIVE; digit2<=NINE; digit3<=THREE; end
      16'd3956: begin digit0<=SIX; digit1<=FIVE; digit2<=NINE; digit3<=THREE; end
      16'd3957: begin digit0<=SEVEN; digit1<=FIVE; digit2<=NINE; digit3<=THREE; end
      16'd3958: begin digit0<=EIGHT; digit1<=FIVE; digit2<=NINE; digit3<=THREE; end
      16'd3959: begin digit0<=NINE; digit1<=FIVE; digit2<=NINE; digit3<=THREE; end
      16'd3960: begin digit0<=ZERO; digit1<=SIX; digit2<=NINE; digit3<=THREE; end
      16'd3961: begin digit0<=ONE; digit1<=SIX; digit2<=NINE; digit3<=THREE; end
      16'd3962: begin digit0<=TWO; digit1<=SIX; digit2<=NINE; digit3<=THREE; end
      16'd3963: begin digit0<=THREE; digit1<=SIX; digit2<=NINE; digit3<=THREE; end
      16'd3964: begin digit0<=FOUR; digit1<=SIX; digit2<=NINE; digit3<=THREE; end
      16'd3965: begin digit0<=FIVE; digit1<=SIX; digit2<=NINE; digit3<=THREE; end
      16'd3966: begin digit0<=SIX; digit1<=SIX; digit2<=NINE; digit3<=THREE; end
      16'd3967: begin digit0<=SEVEN; digit1<=SIX; digit2<=NINE; digit3<=THREE; end
      16'd3968: begin digit0<=EIGHT; digit1<=SIX; digit2<=NINE; digit3<=THREE; end
      16'd3969: begin digit0<=NINE; digit1<=SIX; digit2<=NINE; digit3<=THREE; end
      16'd3970: begin digit0<=ZERO; digit1<=SEVEN; digit2<=NINE; digit3<=THREE; end
      16'd3971: begin digit0<=ONE; digit1<=SEVEN; digit2<=NINE; digit3<=THREE; end
      16'd3972: begin digit0<=TWO; digit1<=SEVEN; digit2<=NINE; digit3<=THREE; end
      16'd3973: begin digit0<=THREE; digit1<=SEVEN; digit2<=NINE; digit3<=THREE; end
      16'd3974: begin digit0<=FOUR; digit1<=SEVEN; digit2<=NINE; digit3<=THREE; end
      16'd3975: begin digit0<=FIVE; digit1<=SEVEN; digit2<=NINE; digit3<=THREE; end
      16'd3976: begin digit0<=SIX; digit1<=SEVEN; digit2<=NINE; digit3<=THREE; end
      16'd3977: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=NINE; digit3<=THREE; end
      16'd3978: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=NINE; digit3<=THREE; end
      16'd3979: begin digit0<=NINE; digit1<=SEVEN; digit2<=NINE; digit3<=THREE; end
      16'd3980: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=THREE; end
      16'd3981: begin digit0<=ONE; digit1<=EIGHT; digit2<=NINE; digit3<=THREE; end
      16'd3982: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=THREE; end
      16'd3983: begin digit0<=THREE; digit1<=EIGHT; digit2<=NINE; digit3<=THREE; end
      16'd3984: begin digit0<=FOUR; digit1<=EIGHT; digit2<=NINE; digit3<=THREE; end
      16'd3985: begin digit0<=FIVE; digit1<=EIGHT; digit2<=NINE; digit3<=THREE; end
      16'd3986: begin digit0<=SIX; digit1<=EIGHT; digit2<=NINE; digit3<=THREE; end
      16'd3987: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=NINE; digit3<=THREE; end
      16'd3988: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=NINE; digit3<=THREE; end
      16'd3989: begin digit0<=NINE; digit1<=EIGHT; digit2<=NINE; digit3<=THREE; end
      16'd3990: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=THREE; end
      16'd3991: begin digit0<=ONE; digit1<=NINE; digit2<=NINE; digit3<=THREE; end
      16'd3992: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=THREE; end
      16'd3993: begin digit0<=THREE; digit1<=NINE; digit2<=NINE; digit3<=THREE; end
      16'd3994: begin digit0<=FOUR; digit1<=NINE; digit2<=NINE; digit3<=THREE; end
      16'd3995: begin digit0<=FIVE; digit1<=NINE; digit2<=NINE; digit3<=THREE; end
      16'd3996: begin digit0<=SIX; digit1<=NINE; digit2<=NINE; digit3<=THREE; end
      16'd3997: begin digit0<=SEVEN; digit1<=NINE; digit2<=NINE; digit3<=THREE; end
      16'd3998: begin digit0<=EIGHT; digit1<=NINE; digit2<=NINE; digit3<=THREE; end
      16'd3999: begin digit0<=NINE; digit1<=NINE; digit2<=NINE; digit3<=THREE; end
	  16'd4000: begin digit0<=ZERO; digit1<=ZERO; digit2<=ZERO; digit3<=FOUR; end
      16'd4001: begin digit0<=ONE; digit1<=ZERO; digit2<=ZERO; digit3<=FOUR; end
      16'd4002: begin digit0<=TWO; digit1<=ZERO; digit2<=ZERO; digit3<=FOUR; end
      16'd4003: begin digit0<=THREE; digit1<=ZERO; digit2<=ZERO; digit3<=FOUR; end
      16'd4004: begin digit0<=FOUR; digit1<=ZERO; digit2<=ZERO; digit3<=FOUR; end
      16'd4005: begin digit0<=FIVE; digit1<=ZERO; digit2<=ZERO; digit3<=FOUR; end
      16'd4006: begin digit0<=SIX; digit1<=ZERO; digit2<=ZERO; digit3<=FOUR; end
      16'd4007: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ZERO; digit3<=FOUR; end
      16'd4008: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ZERO; digit3<=FOUR; end
      16'd4009: begin digit0<=NINE; digit1<=ZERO; digit2<=ZERO; digit3<=FOUR; end
      16'd4010: begin digit0<=ZERO; digit1<=ONE; digit2<=ZERO; digit3<=FOUR; end
      16'd4011: begin digit0<=ONE; digit1<=ONE; digit2<=ZERO; digit3<=FOUR; end
      16'd4012: begin digit0<=TWO; digit1<=ONE; digit2<=ZERO; digit3<=FOUR; end
      16'd4013: begin digit0<=THREE; digit1<=ONE; digit2<=ZERO; digit3<=FOUR; end
      16'd4014: begin digit0<=FOUR; digit1<=ONE; digit2<=ZERO; digit3<=FOUR; end
      16'd4015: begin digit0<=FIVE; digit1<=ONE; digit2<=ZERO; digit3<=FOUR; end
      16'd4016: begin digit0<=SIX; digit1<=ONE; digit2<=ZERO; digit3<=FOUR; end
      16'd4017: begin digit0<=SEVEN; digit1<=ONE; digit2<=ZERO; digit3<=FOUR; end
      16'd4018: begin digit0<=EIGHT; digit1<=ONE; digit2<=ZERO; digit3<=FOUR; end
      16'd4019: begin digit0<=NINE; digit1<=ONE; digit2<=ZERO; digit3<=FOUR; end
      16'd4020: begin digit0<=ZERO; digit1<=TWO; digit2<=ZERO; digit3<=FOUR; end
      16'd4021: begin digit0<=ONE; digit1<=TWO; digit2<=ZERO; digit3<=FOUR; end
      16'd4022: begin digit0<=TWO; digit1<=TWO; digit2<=ZERO; digit3<=FOUR; end
      16'd4023: begin digit0<=THREE; digit1<=TWO; digit2<=ZERO; digit3<=FOUR; end
      16'd4024: begin digit0<=FOUR; digit1<=TWO; digit2<=ZERO; digit3<=FOUR; end
      16'd4025: begin digit0<=FIVE; digit1<=TWO; digit2<=ZERO; digit3<=FOUR; end
      16'd4026: begin digit0<=SIX; digit1<=TWO; digit2<=ZERO; digit3<=FOUR; end
      16'd4027: begin digit0<=SEVEN; digit1<=TWO; digit2<=ZERO; digit3<=FOUR; end
      16'd4028: begin digit0<=EIGHT; digit1<=TWO; digit2<=ZERO; digit3<=FOUR; end
      16'd4029: begin digit0<=NINE; digit1<=TWO; digit2<=ZERO; digit3<=FOUR; end
      16'd4030: begin digit0<=ZERO; digit1<=THREE; digit2<=ZERO; digit3<=FOUR; end
      16'd4031: begin digit0<=ONE; digit1<=THREE; digit2<=ZERO; digit3<=FOUR; end
      16'd4032: begin digit0<=TWO; digit1<=THREE; digit2<=ZERO; digit3<=FOUR; end
      16'd4033: begin digit0<=THREE; digit1<=THREE; digit2<=ZERO; digit3<=FOUR; end
      16'd4034: begin digit0<=FOUR; digit1<=THREE; digit2<=ZERO; digit3<=FOUR; end
      16'd4035: begin digit0<=FIVE; digit1<=THREE; digit2<=ZERO; digit3<=FOUR; end
      16'd4036: begin digit0<=SIX; digit1<=THREE; digit2<=ZERO; digit3<=FOUR; end
      16'd4037: begin digit0<=SEVEN; digit1<=THREE; digit2<=ZERO; digit3<=FOUR; end
      16'd4038: begin digit0<=EIGHT; digit1<=THREE; digit2<=ZERO; digit3<=FOUR; end
      16'd4039: begin digit0<=NINE; digit1<=THREE; digit2<=ZERO; digit3<=FOUR; end
      16'd4040: begin digit0<=ZERO; digit1<=FOUR; digit2<=ZERO; digit3<=FOUR; end
      16'd4041: begin digit0<=ONE; digit1<=FOUR; digit2<=ZERO; digit3<=FOUR; end
      16'd4042: begin digit0<=TWO; digit1<=FOUR; digit2<=ZERO; digit3<=FOUR; end
      16'd4043: begin digit0<=THREE; digit1<=FOUR; digit2<=ZERO; digit3<=FOUR; end
      16'd4044: begin digit0<=FOUR; digit1<=FOUR; digit2<=ZERO; digit3<=FOUR; end
      16'd4045: begin digit0<=FIVE; digit1<=FOUR; digit2<=ZERO; digit3<=FOUR; end
      16'd4046: begin digit0<=SIX; digit1<=FOUR; digit2<=ZERO; digit3<=FOUR; end
      16'd4047: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ZERO; digit3<=FOUR; end
      16'd4048: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ZERO; digit3<=FOUR; end
      16'd4049: begin digit0<=NINE; digit1<=FOUR; digit2<=ZERO; digit3<=FOUR; end
      16'd4050: begin digit0<=ZERO; digit1<=FIVE; digit2<=ZERO; digit3<=FOUR; end
      16'd4051: begin digit0<=ONE; digit1<=FIVE; digit2<=ZERO; digit3<=FOUR; end
      16'd4052: begin digit0<=TWO; digit1<=FIVE; digit2<=ZERO; digit3<=FOUR; end
      16'd4053: begin digit0<=THREE; digit1<=FIVE; digit2<=ZERO; digit3<=FOUR; end
      16'd4054: begin digit0<=FOUR; digit1<=FIVE; digit2<=ZERO; digit3<=FOUR; end
      16'd4055: begin digit0<=FIVE; digit1<=FIVE; digit2<=ZERO; digit3<=FOUR; end
      16'd4056: begin digit0<=SIX; digit1<=FIVE; digit2<=ZERO; digit3<=FOUR; end
      16'd4057: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ZERO; digit3<=FOUR; end
      16'd4058: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ZERO; digit3<=FOUR; end
      16'd4059: begin digit0<=NINE; digit1<=FIVE; digit2<=ZERO; digit3<=FOUR; end
      16'd4060: begin digit0<=ZERO; digit1<=SIX; digit2<=ZERO; digit3<=FOUR; end
      16'd4061: begin digit0<=ONE; digit1<=SIX; digit2<=ZERO; digit3<=FOUR; end
      16'd4062: begin digit0<=TWO; digit1<=SIX; digit2<=ZERO; digit3<=FOUR; end
      16'd4063: begin digit0<=THREE; digit1<=SIX; digit2<=ZERO; digit3<=FOUR; end
      16'd4064: begin digit0<=FOUR; digit1<=SIX; digit2<=ZERO; digit3<=FOUR; end
      16'd4065: begin digit0<=FIVE; digit1<=SIX; digit2<=ZERO; digit3<=FOUR; end
      16'd4066: begin digit0<=SIX; digit1<=SIX; digit2<=ZERO; digit3<=FOUR; end
      16'd4067: begin digit0<=SEVEN; digit1<=SIX; digit2<=ZERO; digit3<=FOUR; end
      16'd4068: begin digit0<=EIGHT; digit1<=SIX; digit2<=ZERO; digit3<=FOUR; end
      16'd4069: begin digit0<=NINE; digit1<=SIX; digit2<=ZERO; digit3<=FOUR; end
      16'd4070: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ZERO; digit3<=FOUR; end
      16'd4071: begin digit0<=ONE; digit1<=SEVEN; digit2<=ZERO; digit3<=FOUR; end
      16'd4072: begin digit0<=TWO; digit1<=SEVEN; digit2<=ZERO; digit3<=FOUR; end
      16'd4073: begin digit0<=THREE; digit1<=SEVEN; digit2<=ZERO; digit3<=FOUR; end
      16'd4074: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ZERO; digit3<=FOUR; end
      16'd4075: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ZERO; digit3<=FOUR; end
      16'd4076: begin digit0<=SIX; digit1<=SEVEN; digit2<=ZERO; digit3<=FOUR; end
      16'd4077: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ZERO; digit3<=FOUR; end
      16'd4078: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ZERO; digit3<=FOUR; end
      16'd4079: begin digit0<=NINE; digit1<=SEVEN; digit2<=ZERO; digit3<=FOUR; end
      16'd4080: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ZERO; digit3<=FOUR; end
      16'd4081: begin digit0<=ONE; digit1<=EIGHT; digit2<=ZERO; digit3<=FOUR; end
      16'd4082: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ZERO; digit3<=FOUR; end
      16'd4083: begin digit0<=THREE; digit1<=EIGHT; digit2<=ZERO; digit3<=FOUR; end
      16'd4084: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ZERO; digit3<=FOUR; end
      16'd4085: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ZERO; digit3<=FOUR; end
      16'd4086: begin digit0<=SIX; digit1<=EIGHT; digit2<=ZERO; digit3<=FOUR; end
      16'd4087: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ZERO; digit3<=FOUR; end
      16'd4088: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ZERO; digit3<=FOUR; end
      16'd4089: begin digit0<=NINE; digit1<=EIGHT; digit2<=ZERO; digit3<=FOUR; end
      16'd4090: begin digit0<=ZERO; digit1<=NINE; digit2<=ZERO; digit3<=FOUR; end
      16'd4091: begin digit0<=ONE; digit1<=NINE; digit2<=ZERO; digit3<=FOUR; end
      16'd4092: begin digit0<=ZERO; digit1<=NINE; digit2<=ZERO; digit3<=FOUR; end
      16'd4093: begin digit0<=THREE; digit1<=NINE; digit2<=ZERO; digit3<=FOUR; end
      16'd4094: begin digit0<=FOUR; digit1<=NINE; digit2<=ZERO; digit3<=FOUR; end
      16'd4095: begin digit0<=FIVE; digit1<=NINE; digit2<=ZERO; digit3<=FOUR; end
      16'd4096: begin digit0<=SIX; digit1<=NINE; digit2<=ZERO; digit3<=FOUR; end
      16'd4097: begin digit0<=SEVEN; digit1<=NINE; digit2<=ZERO; digit3<=FOUR; end
      16'd4098: begin digit0<=EIGHT; digit1<=NINE; digit2<=ZERO; digit3<=FOUR; end
      16'd4099: begin digit0<=NINE; digit1<=NINE; digit2<=ZERO; digit3<=FOUR; end
	  16'd4100: begin digit0<=ZERO; digit1<=ZERO; digit2<=ONE; digit3<=FOUR; end
      16'd4101: begin digit0<=ONE; digit1<=ZERO; digit2<=ONE; digit3<=FOUR; end
      16'd4102: begin digit0<=TWO; digit1<=ZERO; digit2<=ONE; digit3<=FOUR; end
      16'd4103: begin digit0<=THREE; digit1<=ZERO; digit2<=ONE; digit3<=FOUR; end
      16'd4104: begin digit0<=FOUR; digit1<=ZERO; digit2<=ONE; digit3<=FOUR; end
      16'd4105: begin digit0<=FIVE; digit1<=ZERO; digit2<=ONE; digit3<=FOUR; end
      16'd4106: begin digit0<=SIX; digit1<=ZERO; digit2<=ONE; digit3<=FOUR; end
      16'd4107: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ONE; digit3<=FOUR; end
      16'd4108: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ONE; digit3<=FOUR; end
      16'd4109: begin digit0<=NINE; digit1<=ZERO; digit2<=ONE; digit3<=FOUR; end
      16'd4110: begin digit0<=ZERO; digit1<=ONE; digit2<=ONE; digit3<=FOUR; end
      16'd4111: begin digit0<=ONE; digit1<=ONE; digit2<=ONE; digit3<=FOUR; end
      16'd4112: begin digit0<=TWO; digit1<=ONE; digit2<=ONE; digit3<=FOUR; end
      16'd4113: begin digit0<=THREE; digit1<=ONE; digit2<=ONE; digit3<=FOUR; end
      16'd4114: begin digit0<=FOUR; digit1<=ONE; digit2<=ONE; digit3<=FOUR; end
      16'd4115: begin digit0<=FIVE; digit1<=ONE; digit2<=ONE; digit3<=FOUR; end
      16'd4116: begin digit0<=SIX; digit1<=ONE; digit2<=ONE; digit3<=FOUR; end
      16'd4117: begin digit0<=SEVEN; digit1<=ONE; digit2<=ONE; digit3<=FOUR; end
      16'd4118: begin digit0<=EIGHT; digit1<=ONE; digit2<=ONE; digit3<=FOUR; end
      16'd4119: begin digit0<=NINE; digit1<=ONE; digit2<=ONE; digit3<=FOUR; end
      16'd4120: begin digit0<=ZERO; digit1<=TWO; digit2<=ONE; digit3<=FOUR; end
      16'd4121: begin digit0<=ONE; digit1<=TWO; digit2<=ONE; digit3<=FOUR; end
      16'd4122: begin digit0<=TWO; digit1<=TWO; digit2<=ONE; digit3<=FOUR; end
      16'd4123: begin digit0<=THREE; digit1<=TWO; digit2<=ONE; digit3<=FOUR; end
      16'd4124: begin digit0<=FOUR; digit1<=TWO; digit2<=ONE; digit3<=FOUR; end
      16'd4125: begin digit0<=FIVE; digit1<=TWO; digit2<=ONE; digit3<=FOUR; end
      16'd4126: begin digit0<=SIX; digit1<=TWO; digit2<=ONE; digit3<=FOUR; end
      16'd4127: begin digit0<=SEVEN; digit1<=TWO; digit2<=ONE; digit3<=FOUR; end
      16'd4128: begin digit0<=EIGHT; digit1<=TWO; digit2<=ONE; digit3<=FOUR; end
      16'd4129: begin digit0<=NINE; digit1<=TWO; digit2<=ONE; digit3<=FOUR; end
      16'd4130: begin digit0<=ZERO; digit1<=THREE; digit2<=ONE; digit3<=FOUR; end
      16'd4131: begin digit0<=ONE; digit1<=THREE; digit2<=ONE; digit3<=FOUR; end
      16'd4132: begin digit0<=TWO; digit1<=THREE; digit2<=ONE; digit3<=FOUR; end
      16'd4133: begin digit0<=THREE; digit1<=THREE; digit2<=ONE; digit3<=FOUR; end
      16'd4134: begin digit0<=FOUR; digit1<=THREE; digit2<=ONE; digit3<=FOUR; end
      16'd4135: begin digit0<=FIVE; digit1<=THREE; digit2<=ONE; digit3<=FOUR; end
      16'd4136: begin digit0<=SIX; digit1<=THREE; digit2<=ONE; digit3<=FOUR; end
      16'd4137: begin digit0<=SEVEN; digit1<=THREE; digit2<=ONE; digit3<=FOUR; end
      16'd4138: begin digit0<=EIGHT; digit1<=THREE; digit2<=ONE; digit3<=FOUR; end
      16'd4139: begin digit0<=NINE; digit1<=THREE; digit2<=ONE; digit3<=FOUR; end
      16'd4140: begin digit0<=ZERO; digit1<=FOUR; digit2<=ONE; digit3<=FOUR; end
      16'd4141: begin digit0<=ONE; digit1<=FOUR; digit2<=ONE; digit3<=FOUR; end
      16'd4142: begin digit0<=TWO; digit1<=FOUR; digit2<=ONE; digit3<=FOUR; end
      16'd4143: begin digit0<=THREE; digit1<=FOUR; digit2<=ONE; digit3<=FOUR; end
      16'd4144: begin digit0<=FOUR; digit1<=FOUR; digit2<=ONE; digit3<=FOUR; end
      16'd4145: begin digit0<=FIVE; digit1<=FOUR; digit2<=ONE; digit3<=FOUR; end
      16'd4146: begin digit0<=SIX; digit1<=FOUR; digit2<=ONE; digit3<=FOUR; end
      16'd4147: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ONE; digit3<=FOUR; end
      16'd4148: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ONE; digit3<=FOUR; end
      16'd4149: begin digit0<=NINE; digit1<=FOUR; digit2<=ONE; digit3<=FOUR; end
      16'd4150: begin digit0<=ZERO; digit1<=FIVE; digit2<=ONE; digit3<=FOUR; end
      16'd4151: begin digit0<=ONE; digit1<=FIVE; digit2<=ONE; digit3<=FOUR; end
      16'd4152: begin digit0<=TWO; digit1<=FIVE; digit2<=ONE; digit3<=FOUR; end
      16'd4153: begin digit0<=THREE; digit1<=FIVE; digit2<=ONE; digit3<=FOUR; end
      16'd4154: begin digit0<=FOUR; digit1<=FIVE; digit2<=ONE; digit3<=FOUR; end
      16'd4155: begin digit0<=FIVE; digit1<=FIVE; digit2<=ONE; digit3<=FOUR; end
      16'd4156: begin digit0<=SIX; digit1<=FIVE; digit2<=ONE; digit3<=FOUR; end
      16'd4157: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ONE; digit3<=FOUR; end
      16'd4158: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ONE; digit3<=FOUR; end
      16'd4159: begin digit0<=NINE; digit1<=FIVE; digit2<=ONE; digit3<=FOUR; end
      16'd4160: begin digit0<=ZERO; digit1<=SIX; digit2<=ONE; digit3<=FOUR; end
      16'd4161: begin digit0<=ONE; digit1<=SIX; digit2<=ONE; digit3<=FOUR; end
      16'd4162: begin digit0<=TWO; digit1<=SIX; digit2<=ONE; digit3<=FOUR; end
      16'd4163: begin digit0<=THREE; digit1<=SIX; digit2<=ONE; digit3<=FOUR; end
      16'd4164: begin digit0<=FOUR; digit1<=SIX; digit2<=ONE; digit3<=FOUR; end
      16'd4165: begin digit0<=FIVE; digit1<=SIX; digit2<=ONE; digit3<=FOUR; end
      16'd4166: begin digit0<=SIX; digit1<=SIX; digit2<=ONE; digit3<=FOUR; end
      16'd4167: begin digit0<=SEVEN; digit1<=SIX; digit2<=ONE; digit3<=FOUR; end
      16'd4168: begin digit0<=EIGHT; digit1<=SIX; digit2<=ONE; digit3<=FOUR; end
      16'd4169: begin digit0<=NINE; digit1<=SIX; digit2<=ONE; digit3<=FOUR; end
      16'd4170: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ONE; digit3<=FOUR; end
      16'd4171: begin digit0<=ONE; digit1<=SEVEN; digit2<=ONE; digit3<=FOUR; end
      16'd4172: begin digit0<=TWO; digit1<=SEVEN; digit2<=ONE; digit3<=FOUR; end
      16'd4173: begin digit0<=THREE; digit1<=SEVEN; digit2<=ONE; digit3<=FOUR; end
      16'd4174: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ONE; digit3<=FOUR; end
      16'd4175: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ONE; digit3<=FOUR; end
      16'd4176: begin digit0<=SIX; digit1<=SEVEN; digit2<=ONE; digit3<=FOUR; end
      16'd4177: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ONE; digit3<=FOUR; end
      16'd4178: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ONE; digit3<=FOUR; end
      16'd4179: begin digit0<=NINE; digit1<=SEVEN; digit2<=ONE; digit3<=FOUR; end
      16'd4180: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=FOUR; end
      16'd4181: begin digit0<=ONE; digit1<=EIGHT; digit2<=ONE; digit3<=FOUR; end
      16'd4182: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=FOUR; end
      16'd4183: begin digit0<=THREE; digit1<=EIGHT; digit2<=ONE; digit3<=FOUR; end
      16'd4184: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ONE; digit3<=FOUR; end
      16'd4185: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ONE; digit3<=FOUR; end
      16'd4186: begin digit0<=SIX; digit1<=EIGHT; digit2<=ONE; digit3<=FOUR; end
      16'd4187: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ONE; digit3<=FOUR; end
      16'd4188: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ONE; digit3<=FOUR; end
      16'd4189: begin digit0<=NINE; digit1<=EIGHT; digit2<=ONE; digit3<=FOUR; end
      16'd4190: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=FOUR; end
      16'd4191: begin digit0<=ONE; digit1<=NINE; digit2<=ONE; digit3<=FOUR; end
      16'd4192: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=FOUR; end
      16'd4193: begin digit0<=THREE; digit1<=NINE; digit2<=ONE; digit3<=FOUR; end
      16'd4194: begin digit0<=FOUR; digit1<=NINE; digit2<=ONE; digit3<=FOUR; end
      16'd4195: begin digit0<=FIVE; digit1<=NINE; digit2<=ONE; digit3<=FOUR; end
      16'd4196: begin digit0<=SIX; digit1<=NINE; digit2<=ONE; digit3<=FOUR; end
      16'd4197: begin digit0<=SEVEN; digit1<=NINE; digit2<=ONE; digit3<=FOUR; end
      16'd4198: begin digit0<=EIGHT; digit1<=NINE; digit2<=ONE; digit3<=FOUR; end
      16'd4199: begin digit0<=NINE; digit1<=NINE; digit2<=ONE; digit3<=FOUR; end
	  16'd4200: begin digit0<=ZERO; digit1<=ZERO; digit2<=TWO; digit3<=FOUR; end
      16'd4201: begin digit0<=ONE; digit1<=ZERO; digit2<=TWO; digit3<=FOUR; end
      16'd4202: begin digit0<=TWO; digit1<=ZERO; digit2<=TWO; digit3<=FOUR; end
      16'd4203: begin digit0<=THREE; digit1<=ZERO; digit2<=TWO; digit3<=FOUR; end
      16'd4204: begin digit0<=FOUR; digit1<=ZERO; digit2<=TWO; digit3<=FOUR; end
      16'd4205: begin digit0<=FIVE; digit1<=ZERO; digit2<=TWO; digit3<=FOUR; end
      16'd4206: begin digit0<=SIX; digit1<=ZERO; digit2<=TWO; digit3<=FOUR; end
      16'd4207: begin digit0<=SEVEN; digit1<=ZERO; digit2<=TWO; digit3<=FOUR; end
      16'd4208: begin digit0<=EIGHT; digit1<=ZERO; digit2<=TWO; digit3<=FOUR; end
      16'd4209: begin digit0<=NINE; digit1<=ZERO; digit2<=TWO; digit3<=FOUR; end
      16'd4210: begin digit0<=ZERO; digit1<=ONE; digit2<=TWO; digit3<=FOUR; end
      16'd4211: begin digit0<=ONE; digit1<=ONE; digit2<=TWO; digit3<=FOUR; end
      16'd4212: begin digit0<=TWO; digit1<=ONE; digit2<=TWO; digit3<=FOUR; end
      16'd4213: begin digit0<=THREE; digit1<=ONE; digit2<=TWO; digit3<=FOUR; end
      16'd4214: begin digit0<=FOUR; digit1<=ONE; digit2<=TWO; digit3<=FOUR; end
      16'd4215: begin digit0<=FIVE; digit1<=ONE; digit2<=TWO; digit3<=FOUR; end
      16'd4216: begin digit0<=SIX; digit1<=ONE; digit2<=TWO; digit3<=FOUR; end
      16'd4217: begin digit0<=SEVEN; digit1<=ONE; digit2<=TWO; digit3<=FOUR; end
      16'd4218: begin digit0<=EIGHT; digit1<=ONE; digit2<=TWO; digit3<=FOUR; end
      16'd4219: begin digit0<=NINE; digit1<=ONE; digit2<=TWO; digit3<=FOUR; end
      16'd4220: begin digit0<=ZERO; digit1<=TWO; digit2<=TWO; digit3<=FOUR; end
      16'd4221: begin digit0<=ONE; digit1<=TWO; digit2<=TWO; digit3<=FOUR; end
      16'd4222: begin digit0<=TWO; digit1<=TWO; digit2<=TWO; digit3<=FOUR; end
      16'd4223: begin digit0<=THREE; digit1<=TWO; digit2<=TWO; digit3<=FOUR; end
      16'd4224: begin digit0<=FOUR; digit1<=TWO; digit2<=TWO; digit3<=FOUR; end
      16'd4225: begin digit0<=FIVE; digit1<=TWO; digit2<=TWO; digit3<=FOUR; end
      16'd4226: begin digit0<=SIX; digit1<=TWO; digit2<=TWO; digit3<=FOUR; end
      16'd4227: begin digit0<=SEVEN; digit1<=TWO; digit2<=TWO; digit3<=FOUR; end
      16'd4228: begin digit0<=EIGHT; digit1<=TWO; digit2<=TWO; digit3<=FOUR; end
      16'd4229: begin digit0<=NINE; digit1<=TWO; digit2<=TWO; digit3<=FOUR; end
      16'd4230: begin digit0<=ZERO; digit1<=THREE; digit2<=TWO; digit3<=FOUR; end
      16'd4231: begin digit0<=ONE; digit1<=THREE; digit2<=TWO; digit3<=FOUR; end
      16'd4232: begin digit0<=TWO; digit1<=THREE; digit2<=TWO; digit3<=FOUR; end
      16'd4233: begin digit0<=THREE; digit1<=THREE; digit2<=TWO; digit3<=FOUR; end
      16'd4234: begin digit0<=FOUR; digit1<=THREE; digit2<=TWO; digit3<=FOUR; end
      16'd4235: begin digit0<=FIVE; digit1<=THREE; digit2<=TWO; digit3<=FOUR; end
      16'd4236: begin digit0<=SIX; digit1<=THREE; digit2<=TWO; digit3<=FOUR; end
      16'd4237: begin digit0<=SEVEN; digit1<=THREE; digit2<=TWO; digit3<=FOUR; end
      16'd4238: begin digit0<=EIGHT; digit1<=THREE; digit2<=TWO; digit3<=FOUR; end
      16'd4239: begin digit0<=NINE; digit1<=THREE; digit2<=TWO; digit3<=FOUR; end
      16'd4240: begin digit0<=ZERO; digit1<=FOUR; digit2<=TWO; digit3<=FOUR; end
      16'd4241: begin digit0<=ONE; digit1<=FOUR; digit2<=TWO; digit3<=FOUR; end
      16'd4242: begin digit0<=TWO; digit1<=FOUR; digit2<=TWO; digit3<=FOUR; end
      16'd4243: begin digit0<=THREE; digit1<=FOUR; digit2<=TWO; digit3<=FOUR; end
      16'd4244: begin digit0<=FOUR; digit1<=FOUR; digit2<=TWO; digit3<=FOUR; end
      16'd4245: begin digit0<=FIVE; digit1<=FOUR; digit2<=TWO; digit3<=FOUR; end
      16'd4246: begin digit0<=SIX; digit1<=FOUR; digit2<=TWO; digit3<=FOUR; end
      16'd4247: begin digit0<=SEVEN; digit1<=FOUR; digit2<=TWO; digit3<=FOUR; end
      16'd4248: begin digit0<=EIGHT; digit1<=FOUR; digit2<=TWO; digit3<=FOUR; end
      16'd4249: begin digit0<=NINE; digit1<=FOUR; digit2<=TWO; digit3<=FOUR; end
      16'd4250: begin digit0<=ZERO; digit1<=FIVE; digit2<=TWO; digit3<=FOUR; end
      16'd4251: begin digit0<=ONE; digit1<=FIVE; digit2<=TWO; digit3<=FOUR; end
      16'd4252: begin digit0<=TWO; digit1<=FIVE; digit2<=TWO; digit3<=FOUR; end
      16'd4253: begin digit0<=THREE; digit1<=FIVE; digit2<=TWO; digit3<=FOUR; end
      16'd4254: begin digit0<=FOUR; digit1<=FIVE; digit2<=TWO; digit3<=FOUR; end
      16'd4255: begin digit0<=FIVE; digit1<=FIVE; digit2<=TWO; digit3<=FOUR; end
      16'd4256: begin digit0<=SIX; digit1<=FIVE; digit2<=TWO; digit3<=FOUR; end
      16'd4257: begin digit0<=SEVEN; digit1<=FIVE; digit2<=TWO; digit3<=FOUR; end
      16'd4258: begin digit0<=EIGHT; digit1<=FIVE; digit2<=TWO; digit3<=FOUR; end
      16'd4259: begin digit0<=NINE; digit1<=FIVE; digit2<=TWO; digit3<=FOUR; end
      16'd4260: begin digit0<=ZERO; digit1<=SIX; digit2<=TWO; digit3<=FOUR; end
      16'd4261: begin digit0<=ONE; digit1<=SIX; digit2<=TWO; digit3<=FOUR; end
      16'd4262: begin digit0<=TWO; digit1<=SIX; digit2<=TWO; digit3<=FOUR; end
      16'd4263: begin digit0<=THREE; digit1<=SIX; digit2<=TWO; digit3<=FOUR; end
      16'd4264: begin digit0<=FOUR; digit1<=SIX; digit2<=TWO; digit3<=FOUR; end
      16'd4265: begin digit0<=FIVE; digit1<=SIX; digit2<=TWO; digit3<=FOUR; end
      16'd4266: begin digit0<=SIX; digit1<=SIX; digit2<=TWO; digit3<=FOUR; end
      16'd4267: begin digit0<=SEVEN; digit1<=SIX; digit2<=TWO; digit3<=FOUR; end
      16'd4268: begin digit0<=EIGHT; digit1<=SIX; digit2<=TWO; digit3<=FOUR; end
      16'd4269: begin digit0<=NINE; digit1<=SIX; digit2<=TWO; digit3<=FOUR; end
      16'd4270: begin digit0<=ZERO; digit1<=SEVEN; digit2<=TWO; digit3<=FOUR; end
      16'd4271: begin digit0<=ONE; digit1<=SEVEN; digit2<=TWO; digit3<=FOUR; end
      16'd4272: begin digit0<=TWO; digit1<=SEVEN; digit2<=TWO; digit3<=FOUR; end
      16'd4273: begin digit0<=THREE; digit1<=SEVEN; digit2<=TWO; digit3<=FOUR; end
      16'd4274: begin digit0<=FOUR; digit1<=SEVEN; digit2<=TWO; digit3<=FOUR; end
      16'd4275: begin digit0<=FIVE; digit1<=SEVEN; digit2<=TWO; digit3<=FOUR; end
      16'd4276: begin digit0<=SIX; digit1<=SEVEN; digit2<=TWO; digit3<=FOUR; end
      16'd4277: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=TWO; digit3<=FOUR; end
      16'd4278: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=TWO; digit3<=FOUR; end
      16'd4279: begin digit0<=NINE; digit1<=SEVEN; digit2<=TWO; digit3<=FOUR; end
      16'd4280: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=FOUR; end
      16'd4281: begin digit0<=ONE; digit1<=EIGHT; digit2<=TWO; digit3<=FOUR; end
      16'd4282: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=FOUR; end
      16'd4283: begin digit0<=THREE; digit1<=EIGHT; digit2<=TWO; digit3<=FOUR; end
      16'd4284: begin digit0<=FOUR; digit1<=EIGHT; digit2<=TWO; digit3<=FOUR; end
      16'd4285: begin digit0<=FIVE; digit1<=EIGHT; digit2<=TWO; digit3<=FOUR; end
      16'd4286: begin digit0<=SIX; digit1<=EIGHT; digit2<=TWO; digit3<=FOUR; end
      16'd4287: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=TWO; digit3<=FOUR; end
      16'd4288: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=TWO; digit3<=FOUR; end
      16'd4289: begin digit0<=NINE; digit1<=EIGHT; digit2<=TWO; digit3<=FOUR; end
      16'd4290: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=FOUR; end
      16'd4291: begin digit0<=ONE; digit1<=NINE; digit2<=TWO; digit3<=FOUR; end
      16'd4292: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=FOUR; end
      16'd4293: begin digit0<=THREE; digit1<=NINE; digit2<=TWO; digit3<=FOUR; end
      16'd4294: begin digit0<=FOUR; digit1<=NINE; digit2<=TWO; digit3<=FOUR; end
      16'd4295: begin digit0<=FIVE; digit1<=NINE; digit2<=TWO; digit3<=FOUR; end
      16'd4296: begin digit0<=SIX; digit1<=NINE; digit2<=TWO; digit3<=FOUR; end
      16'd4297: begin digit0<=SEVEN; digit1<=NINE; digit2<=TWO; digit3<=FOUR; end
      16'd4298: begin digit0<=EIGHT; digit1<=NINE; digit2<=TWO; digit3<=FOUR; end
      16'd4299: begin digit0<=NINE; digit1<=NINE; digit2<=TWO; digit3<=FOUR; end
	  16'd4300: begin digit0<=ZERO; digit1<=ZERO; digit2<=THREE; digit3<=FOUR; end
      16'd4301: begin digit0<=ONE; digit1<=ZERO; digit2<=THREE; digit3<=FOUR; end
      16'd4302: begin digit0<=TWO; digit1<=ZERO; digit2<=THREE; digit3<=FOUR; end
      16'd4303: begin digit0<=THREE; digit1<=ZERO; digit2<=THREE; digit3<=FOUR; end
      16'd4304: begin digit0<=FOUR; digit1<=ZERO; digit2<=THREE; digit3<=FOUR; end
      16'd4305: begin digit0<=FIVE; digit1<=ZERO; digit2<=THREE; digit3<=FOUR; end
      16'd4306: begin digit0<=SIX; digit1<=ZERO; digit2<=THREE; digit3<=FOUR; end
      16'd4307: begin digit0<=SEVEN; digit1<=ZERO; digit2<=THREE; digit3<=FOUR; end
      16'd4308: begin digit0<=EIGHT; digit1<=ZERO; digit2<=THREE; digit3<=FOUR; end
      16'd4309: begin digit0<=NINE; digit1<=ZERO; digit2<=THREE; digit3<=FOUR; end
      16'd4310: begin digit0<=ZERO; digit1<=ONE; digit2<=THREE; digit3<=FOUR; end
      16'd4311: begin digit0<=ONE; digit1<=ONE; digit2<=THREE; digit3<=FOUR; end
      16'd4312: begin digit0<=TWO; digit1<=ONE; digit2<=THREE; digit3<=FOUR; end
      16'd4313: begin digit0<=THREE; digit1<=ONE; digit2<=THREE; digit3<=FOUR; end
      16'd4314: begin digit0<=FOUR; digit1<=ONE; digit2<=THREE; digit3<=FOUR; end
      16'd4315: begin digit0<=FIVE; digit1<=ONE; digit2<=THREE; digit3<=FOUR; end
      16'd4316: begin digit0<=SIX; digit1<=ONE; digit2<=THREE; digit3<=FOUR; end
      16'd4317: begin digit0<=SEVEN; digit1<=ONE; digit2<=THREE; digit3<=FOUR; end
      16'd4318: begin digit0<=EIGHT; digit1<=ONE; digit2<=THREE; digit3<=FOUR; end
      16'd4319: begin digit0<=NINE; digit1<=ONE; digit2<=THREE; digit3<=FOUR; end
      16'd4320: begin digit0<=ZERO; digit1<=TWO; digit2<=THREE; digit3<=FOUR; end
      16'd4321: begin digit0<=ONE; digit1<=TWO; digit2<=THREE; digit3<=FOUR; end
      16'd4322: begin digit0<=TWO; digit1<=TWO; digit2<=THREE; digit3<=FOUR; end
      16'd4323: begin digit0<=THREE; digit1<=TWO; digit2<=THREE; digit3<=FOUR; end
      16'd4324: begin digit0<=FOUR; digit1<=TWO; digit2<=THREE; digit3<=FOUR; end
      16'd4325: begin digit0<=FIVE; digit1<=TWO; digit2<=THREE; digit3<=FOUR; end
      16'd4326: begin digit0<=SIX; digit1<=TWO; digit2<=THREE; digit3<=FOUR; end
      16'd4327: begin digit0<=SEVEN; digit1<=TWO; digit2<=THREE; digit3<=FOUR; end
      16'd4328: begin digit0<=EIGHT; digit1<=TWO; digit2<=THREE; digit3<=FOUR; end
      16'd4329: begin digit0<=NINE; digit1<=TWO; digit2<=THREE; digit3<=FOUR; end
      16'd4330: begin digit0<=ZERO; digit1<=THREE; digit2<=THREE; digit3<=FOUR; end
      16'd4331: begin digit0<=ONE; digit1<=THREE; digit2<=THREE; digit3<=FOUR; end
      16'd4332: begin digit0<=TWO; digit1<=THREE; digit2<=THREE; digit3<=FOUR; end
      16'd4333: begin digit0<=THREE; digit1<=THREE; digit2<=THREE; digit3<=FOUR; end
      16'd4334: begin digit0<=FOUR; digit1<=THREE; digit2<=THREE; digit3<=FOUR; end
      16'd4335: begin digit0<=FIVE; digit1<=THREE; digit2<=THREE; digit3<=FOUR; end
      16'd4336: begin digit0<=SIX; digit1<=THREE; digit2<=THREE; digit3<=FOUR; end
      16'd4337: begin digit0<=SEVEN; digit1<=THREE; digit2<=THREE; digit3<=FOUR; end
      16'd4338: begin digit0<=EIGHT; digit1<=THREE; digit2<=THREE; digit3<=FOUR; end
      16'd4339: begin digit0<=NINE; digit1<=THREE; digit2<=THREE; digit3<=FOUR; end
      16'd4340: begin digit0<=ZERO; digit1<=FOUR; digit2<=THREE; digit3<=FOUR; end
      16'd4341: begin digit0<=ONE; digit1<=FOUR; digit2<=THREE; digit3<=FOUR; end
      16'd4342: begin digit0<=TWO; digit1<=FOUR; digit2<=THREE; digit3<=FOUR; end
      16'd4343: begin digit0<=THREE; digit1<=FOUR; digit2<=THREE; digit3<=FOUR; end
      16'd4344: begin digit0<=FOUR; digit1<=FOUR; digit2<=THREE; digit3<=FOUR; end
      16'd4345: begin digit0<=FIVE; digit1<=FOUR; digit2<=THREE; digit3<=FOUR; end
      16'd4346: begin digit0<=SIX; digit1<=FOUR; digit2<=THREE; digit3<=FOUR; end
      16'd4347: begin digit0<=SEVEN; digit1<=FOUR; digit2<=THREE; digit3<=FOUR; end
      16'd4348: begin digit0<=EIGHT; digit1<=FOUR; digit2<=THREE; digit3<=FOUR; end
      16'd4349: begin digit0<=NINE; digit1<=FOUR; digit2<=THREE; digit3<=FOUR; end
      16'd4350: begin digit0<=ZERO; digit1<=FIVE; digit2<=THREE; digit3<=FOUR; end
      16'd4351: begin digit0<=ONE; digit1<=FIVE; digit2<=THREE; digit3<=FOUR; end
      16'd4352: begin digit0<=TWO; digit1<=FIVE; digit2<=THREE; digit3<=FOUR; end
      16'd4353: begin digit0<=THREE; digit1<=FIVE; digit2<=THREE; digit3<=FOUR; end
      16'd4354: begin digit0<=FOUR; digit1<=FIVE; digit2<=THREE; digit3<=FOUR; end
      16'd4355: begin digit0<=FIVE; digit1<=FIVE; digit2<=THREE; digit3<=FOUR; end
      16'd4356: begin digit0<=SIX; digit1<=FIVE; digit2<=THREE; digit3<=FOUR; end
      16'd4357: begin digit0<=SEVEN; digit1<=FIVE; digit2<=THREE; digit3<=FOUR; end
      16'd4358: begin digit0<=EIGHT; digit1<=FIVE; digit2<=THREE; digit3<=FOUR; end
      16'd4359: begin digit0<=NINE; digit1<=FIVE; digit2<=THREE; digit3<=FOUR; end
      16'd4360: begin digit0<=ZERO; digit1<=SIX; digit2<=THREE; digit3<=FOUR; end
      16'd4361: begin digit0<=ONE; digit1<=SIX; digit2<=THREE; digit3<=FOUR; end
      16'd4362: begin digit0<=TWO; digit1<=SIX; digit2<=THREE; digit3<=FOUR; end
      16'd4363: begin digit0<=THREE; digit1<=SIX; digit2<=THREE; digit3<=FOUR; end
      16'd4364: begin digit0<=FOUR; digit1<=SIX; digit2<=THREE; digit3<=FOUR; end
      16'd4365: begin digit0<=FIVE; digit1<=SIX; digit2<=THREE; digit3<=FOUR; end
      16'd4366: begin digit0<=SIX; digit1<=SIX; digit2<=THREE; digit3<=FOUR; end
      16'd4367: begin digit0<=SEVEN; digit1<=SIX; digit2<=THREE; digit3<=FOUR; end
      16'd4368: begin digit0<=EIGHT; digit1<=SIX; digit2<=THREE; digit3<=FOUR; end
      16'd4369: begin digit0<=NINE; digit1<=SIX; digit2<=THREE; digit3<=FOUR; end
      16'd4370: begin digit0<=ZERO; digit1<=SEVEN; digit2<=THREE; digit3<=FOUR; end
      16'd4371: begin digit0<=ONE; digit1<=SEVEN; digit2<=THREE; digit3<=FOUR; end
      16'd4372: begin digit0<=TWO; digit1<=SEVEN; digit2<=THREE; digit3<=FOUR; end
      16'd4373: begin digit0<=THREE; digit1<=SEVEN; digit2<=THREE; digit3<=FOUR; end
      16'd4374: begin digit0<=FOUR; digit1<=SEVEN; digit2<=THREE; digit3<=FOUR; end
      16'd4375: begin digit0<=FIVE; digit1<=SEVEN; digit2<=THREE; digit3<=FOUR; end
      16'd4376: begin digit0<=SIX; digit1<=SEVEN; digit2<=THREE; digit3<=FOUR; end
      16'd4377: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=THREE; digit3<=FOUR; end
      16'd4378: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=THREE; digit3<=FOUR; end
      16'd4379: begin digit0<=NINE; digit1<=SEVEN; digit2<=THREE; digit3<=FOUR; end
      16'd4380: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=FOUR; end
      16'd4381: begin digit0<=ONE; digit1<=EIGHT; digit2<=THREE; digit3<=FOUR; end
      16'd4382: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=FOUR; end
      16'd4383: begin digit0<=THREE; digit1<=EIGHT; digit2<=THREE; digit3<=FOUR; end
      16'd4384: begin digit0<=FOUR; digit1<=EIGHT; digit2<=THREE; digit3<=FOUR; end
      16'd4385: begin digit0<=FIVE; digit1<=EIGHT; digit2<=THREE; digit3<=FOUR; end
      16'd4386: begin digit0<=SIX; digit1<=EIGHT; digit2<=THREE; digit3<=FOUR; end
      16'd4387: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=THREE; digit3<=FOUR; end
      16'd4388: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=THREE; digit3<=FOUR; end
      16'd4389: begin digit0<=NINE; digit1<=EIGHT; digit2<=THREE; digit3<=FOUR; end
      16'd4390: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=FOUR; end
      16'd4391: begin digit0<=ONE; digit1<=NINE; digit2<=THREE; digit3<=FOUR; end
      16'd4392: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=FOUR; end
      16'd4393: begin digit0<=THREE; digit1<=NINE; digit2<=THREE; digit3<=FOUR; end
      16'd4394: begin digit0<=FOUR; digit1<=NINE; digit2<=THREE; digit3<=FOUR; end
      16'd4395: begin digit0<=FIVE; digit1<=NINE; digit2<=THREE; digit3<=FOUR; end
      16'd4396: begin digit0<=SIX; digit1<=NINE; digit2<=THREE; digit3<=FOUR; end
      16'd4397: begin digit0<=SEVEN; digit1<=NINE; digit2<=THREE; digit3<=FOUR; end
      16'd4398: begin digit0<=EIGHT; digit1<=NINE; digit2<=THREE; digit3<=FOUR; end
      16'd4399: begin digit0<=NINE; digit1<=NINE; digit2<=THREE; digit3<=FOUR; end
	  16'd4400: begin digit0<=ZERO; digit1<=ZERO; digit2<=FOUR; digit3<=FOUR; end
      16'd4401: begin digit0<=ONE; digit1<=ZERO; digit2<=FOUR; digit3<=FOUR; end
      16'd4402: begin digit0<=TWO; digit1<=ZERO; digit2<=FOUR; digit3<=FOUR; end
      16'd4403: begin digit0<=THREE; digit1<=ZERO; digit2<=FOUR; digit3<=FOUR; end
      16'd4404: begin digit0<=FOUR; digit1<=ZERO; digit2<=FOUR; digit3<=FOUR; end
      16'd4405: begin digit0<=FIVE; digit1<=ZERO; digit2<=FOUR; digit3<=FOUR; end
      16'd4406: begin digit0<=SIX; digit1<=ZERO; digit2<=FOUR; digit3<=FOUR; end
      16'd4407: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FOUR; digit3<=FOUR; end
      16'd4408: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FOUR; digit3<=FOUR; end
      16'd4409: begin digit0<=NINE; digit1<=ZERO; digit2<=FOUR; digit3<=FOUR; end
      16'd4410: begin digit0<=ZERO; digit1<=ONE; digit2<=FOUR; digit3<=FOUR; end
      16'd4411: begin digit0<=ONE; digit1<=ONE; digit2<=FOUR; digit3<=FOUR; end
      16'd4412: begin digit0<=TWO; digit1<=ONE; digit2<=FOUR; digit3<=FOUR; end
      16'd4413: begin digit0<=THREE; digit1<=ONE; digit2<=FOUR; digit3<=FOUR; end
      16'd4414: begin digit0<=FOUR; digit1<=ONE; digit2<=FOUR; digit3<=FOUR; end
      16'd4415: begin digit0<=FIVE; digit1<=ONE; digit2<=FOUR; digit3<=FOUR; end
      16'd4416: begin digit0<=SIX; digit1<=ONE; digit2<=FOUR; digit3<=FOUR; end
      16'd4417: begin digit0<=SEVEN; digit1<=ONE; digit2<=FOUR; digit3<=FOUR; end
      16'd4418: begin digit0<=EIGHT; digit1<=ONE; digit2<=FOUR; digit3<=FOUR; end
      16'd4419: begin digit0<=NINE; digit1<=ONE; digit2<=FOUR; digit3<=FOUR; end
      16'd4420: begin digit0<=ZERO; digit1<=TWO; digit2<=FOUR; digit3<=FOUR; end
      16'd4421: begin digit0<=ONE; digit1<=TWO; digit2<=FOUR; digit3<=FOUR; end
      16'd4422: begin digit0<=TWO; digit1<=TWO; digit2<=FOUR; digit3<=FOUR; end
      16'd4423: begin digit0<=THREE; digit1<=TWO; digit2<=FOUR; digit3<=FOUR; end
      16'd4424: begin digit0<=FOUR; digit1<=TWO; digit2<=FOUR; digit3<=FOUR; end
      16'd4425: begin digit0<=FIVE; digit1<=TWO; digit2<=FOUR; digit3<=FOUR; end
      16'd4426: begin digit0<=SIX; digit1<=TWO; digit2<=FOUR; digit3<=FOUR; end
      16'd4427: begin digit0<=SEVEN; digit1<=TWO; digit2<=FOUR; digit3<=FOUR; end
      16'd4428: begin digit0<=EIGHT; digit1<=TWO; digit2<=FOUR; digit3<=FOUR; end
      16'd4429: begin digit0<=NINE; digit1<=TWO; digit2<=FOUR; digit3<=FOUR; end
      16'd4430: begin digit0<=ZERO; digit1<=THREE; digit2<=FOUR; digit3<=FOUR; end
      16'd4431: begin digit0<=ONE; digit1<=THREE; digit2<=FOUR; digit3<=FOUR; end
      16'd4432: begin digit0<=TWO; digit1<=THREE; digit2<=FOUR; digit3<=FOUR; end
      16'd4433: begin digit0<=THREE; digit1<=THREE; digit2<=FOUR; digit3<=FOUR; end
      16'd4434: begin digit0<=FOUR; digit1<=THREE; digit2<=FOUR; digit3<=FOUR; end
      16'd4435: begin digit0<=FIVE; digit1<=THREE; digit2<=FOUR; digit3<=FOUR; end
      16'd4436: begin digit0<=SIX; digit1<=THREE; digit2<=FOUR; digit3<=FOUR; end
      16'd4437: begin digit0<=SEVEN; digit1<=THREE; digit2<=FOUR; digit3<=FOUR; end
      16'd4438: begin digit0<=EIGHT; digit1<=THREE; digit2<=FOUR; digit3<=FOUR; end
      16'd4439: begin digit0<=NINE; digit1<=THREE; digit2<=FOUR; digit3<=FOUR; end
      16'd4440: begin digit0<=ZERO; digit1<=FOUR; digit2<=FOUR; digit3<=FOUR; end
      16'd4441: begin digit0<=ONE; digit1<=FOUR; digit2<=FOUR; digit3<=FOUR; end
      16'd4442: begin digit0<=TWO; digit1<=FOUR; digit2<=FOUR; digit3<=FOUR; end
      16'd4443: begin digit0<=THREE; digit1<=FOUR; digit2<=FOUR; digit3<=FOUR; end
      16'd4444: begin digit0<=FOUR; digit1<=FOUR; digit2<=FOUR; digit3<=FOUR; end
      16'd4445: begin digit0<=FIVE; digit1<=FOUR; digit2<=FOUR; digit3<=FOUR; end
      16'd4446: begin digit0<=SIX; digit1<=FOUR; digit2<=FOUR; digit3<=FOUR; end
      16'd4447: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FOUR; digit3<=FOUR; end
      16'd4448: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FOUR; digit3<=FOUR; end
      16'd4449: begin digit0<=NINE; digit1<=FOUR; digit2<=FOUR; digit3<=FOUR; end
      16'd4450: begin digit0<=ZERO; digit1<=FIVE; digit2<=FOUR; digit3<=FOUR; end
      16'd4451: begin digit0<=ONE; digit1<=FIVE; digit2<=FOUR; digit3<=FOUR; end
      16'd4452: begin digit0<=TWO; digit1<=FIVE; digit2<=FOUR; digit3<=FOUR; end
      16'd4453: begin digit0<=THREE; digit1<=FIVE; digit2<=FOUR; digit3<=FOUR; end
      16'd4454: begin digit0<=FOUR; digit1<=FIVE; digit2<=FOUR; digit3<=FOUR; end
      16'd4455: begin digit0<=FIVE; digit1<=FIVE; digit2<=FOUR; digit3<=FOUR; end
      16'd4456: begin digit0<=SIX; digit1<=FIVE; digit2<=FOUR; digit3<=FOUR; end
      16'd4457: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FOUR; digit3<=FOUR; end
      16'd4458: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FOUR; digit3<=FOUR; end
      16'd4459: begin digit0<=NINE; digit1<=FIVE; digit2<=FOUR; digit3<=FOUR; end
      16'd4460: begin digit0<=ZERO; digit1<=SIX; digit2<=FOUR; digit3<=FOUR; end
      16'd4461: begin digit0<=ONE; digit1<=SIX; digit2<=FOUR; digit3<=FOUR; end
      16'd4462: begin digit0<=TWO; digit1<=SIX; digit2<=FOUR; digit3<=FOUR; end
      16'd4463: begin digit0<=THREE; digit1<=SIX; digit2<=FOUR; digit3<=FOUR; end
      16'd4464: begin digit0<=FOUR; digit1<=SIX; digit2<=FOUR; digit3<=FOUR; end
      16'd4465: begin digit0<=FIVE; digit1<=SIX; digit2<=FOUR; digit3<=FOUR; end
      16'd4466: begin digit0<=SIX; digit1<=SIX; digit2<=FOUR; digit3<=FOUR; end
      16'd4467: begin digit0<=SEVEN; digit1<=SIX; digit2<=FOUR; digit3<=FOUR; end
      16'd4468: begin digit0<=EIGHT; digit1<=SIX; digit2<=FOUR; digit3<=FOUR; end
      16'd4469: begin digit0<=NINE; digit1<=SIX; digit2<=FOUR; digit3<=FOUR; end
      16'd4470: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FOUR; digit3<=FOUR; end
      16'd4471: begin digit0<=ONE; digit1<=SEVEN; digit2<=FOUR; digit3<=FOUR; end
      16'd4472: begin digit0<=TWO; digit1<=SEVEN; digit2<=FOUR; digit3<=FOUR; end
      16'd4473: begin digit0<=THREE; digit1<=SEVEN; digit2<=FOUR; digit3<=FOUR; end
      16'd4474: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FOUR; digit3<=FOUR; end
      16'd4475: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FOUR; digit3<=FOUR; end
      16'd4476: begin digit0<=SIX; digit1<=SEVEN; digit2<=FOUR; digit3<=FOUR; end
      16'd4477: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FOUR; digit3<=FOUR; end
      16'd4478: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FOUR; digit3<=FOUR; end
      16'd4479: begin digit0<=NINE; digit1<=SEVEN; digit2<=FOUR; digit3<=FOUR; end
      16'd4480: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=FOUR; end
      16'd4481: begin digit0<=ONE; digit1<=EIGHT; digit2<=FOUR; digit3<=FOUR; end
      16'd4482: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=FOUR; end
      16'd4483: begin digit0<=THREE; digit1<=EIGHT; digit2<=FOUR; digit3<=FOUR; end
      16'd4484: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FOUR; digit3<=FOUR; end
      16'd4485: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FOUR; digit3<=FOUR; end
      16'd4486: begin digit0<=SIX; digit1<=EIGHT; digit2<=FOUR; digit3<=FOUR; end
      16'd4487: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FOUR; digit3<=FOUR; end
      16'd4488: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FOUR; digit3<=FOUR; end
      16'd4489: begin digit0<=NINE; digit1<=EIGHT; digit2<=FOUR; digit3<=FOUR; end
      16'd4490: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=FOUR; end
      16'd4491: begin digit0<=ONE; digit1<=NINE; digit2<=FOUR; digit3<=FOUR; end
      16'd4492: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=FOUR; end
      16'd4493: begin digit0<=THREE; digit1<=NINE; digit2<=FOUR; digit3<=FOUR; end
      16'd4494: begin digit0<=FOUR; digit1<=NINE; digit2<=FOUR; digit3<=FOUR; end
      16'd4495: begin digit0<=FIVE; digit1<=NINE; digit2<=FOUR; digit3<=FOUR; end
      16'd4496: begin digit0<=SIX; digit1<=NINE; digit2<=FOUR; digit3<=FOUR; end
      16'd4497: begin digit0<=SEVEN; digit1<=NINE; digit2<=FOUR; digit3<=FOUR; end
      16'd4498: begin digit0<=EIGHT; digit1<=NINE; digit2<=FOUR; digit3<=FOUR; end
      16'd4499: begin digit0<=NINE; digit1<=NINE; digit2<=FOUR; digit3<=FOUR; end
	  16'd4500: begin digit0<=ZERO; digit1<=ZERO; digit2<=FIVE; digit3<=FOUR; end
      16'd4501: begin digit0<=ONE; digit1<=ZERO; digit2<=FIVE; digit3<=FOUR; end
      16'd4502: begin digit0<=TWO; digit1<=ZERO; digit2<=FIVE; digit3<=FOUR; end
      16'd4503: begin digit0<=THREE; digit1<=ZERO; digit2<=FIVE; digit3<=FOUR; end
      16'd4504: begin digit0<=FOUR; digit1<=ZERO; digit2<=FIVE; digit3<=FOUR; end
      16'd4505: begin digit0<=FIVE; digit1<=ZERO; digit2<=FIVE; digit3<=FOUR; end
      16'd4506: begin digit0<=SIX; digit1<=ZERO; digit2<=FIVE; digit3<=FOUR; end
      16'd4507: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FIVE; digit3<=FOUR; end
      16'd4508: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FIVE; digit3<=FOUR; end
      16'd4509: begin digit0<=NINE; digit1<=ZERO; digit2<=FIVE; digit3<=FOUR; end
      16'd4510: begin digit0<=ZERO; digit1<=ONE; digit2<=FIVE; digit3<=FOUR; end
      16'd4511: begin digit0<=ONE; digit1<=ONE; digit2<=FIVE; digit3<=FOUR; end
      16'd4512: begin digit0<=TWO; digit1<=ONE; digit2<=FIVE; digit3<=FOUR; end
      16'd4513: begin digit0<=THREE; digit1<=ONE; digit2<=FIVE; digit3<=FOUR; end
      16'd4514: begin digit0<=FOUR; digit1<=ONE; digit2<=FIVE; digit3<=FOUR; end
      16'd4515: begin digit0<=FIVE; digit1<=ONE; digit2<=FIVE; digit3<=FOUR; end
      16'd4516: begin digit0<=SIX; digit1<=ONE; digit2<=FIVE; digit3<=FOUR; end
      16'd4517: begin digit0<=SEVEN; digit1<=ONE; digit2<=FIVE; digit3<=FOUR; end
      16'd4518: begin digit0<=EIGHT; digit1<=ONE; digit2<=FIVE; digit3<=FOUR; end
      16'd4519: begin digit0<=NINE; digit1<=ONE; digit2<=FIVE; digit3<=FOUR; end
      16'd4520: begin digit0<=ZERO; digit1<=TWO; digit2<=FIVE; digit3<=FOUR; end
      16'd4521: begin digit0<=ONE; digit1<=TWO; digit2<=FIVE; digit3<=FOUR; end
      16'd4522: begin digit0<=TWO; digit1<=TWO; digit2<=FIVE; digit3<=FOUR; end
      16'd4523: begin digit0<=THREE; digit1<=TWO; digit2<=FIVE; digit3<=FOUR; end
      16'd4524: begin digit0<=FOUR; digit1<=TWO; digit2<=FIVE; digit3<=FOUR; end
      16'd4525: begin digit0<=FIVE; digit1<=TWO; digit2<=FIVE; digit3<=FOUR; end
      16'd4526: begin digit0<=SIX; digit1<=TWO; digit2<=FIVE; digit3<=FOUR; end
      16'd4527: begin digit0<=SEVEN; digit1<=TWO; digit2<=FIVE; digit3<=FOUR; end
      16'd4528: begin digit0<=EIGHT; digit1<=TWO; digit2<=FIVE; digit3<=FOUR; end
      16'd4529: begin digit0<=NINE; digit1<=TWO; digit2<=FIVE; digit3<=FOUR; end
      16'd4530: begin digit0<=ZERO; digit1<=THREE; digit2<=FIVE; digit3<=FOUR; end
      16'd4531: begin digit0<=ONE; digit1<=THREE; digit2<=FIVE; digit3<=FOUR; end
      16'd4532: begin digit0<=TWO; digit1<=THREE; digit2<=FIVE; digit3<=FOUR; end
      16'd4533: begin digit0<=THREE; digit1<=THREE; digit2<=FIVE; digit3<=FOUR; end
      16'd4534: begin digit0<=FOUR; digit1<=THREE; digit2<=FIVE; digit3<=FOUR; end
      16'd4535: begin digit0<=FIVE; digit1<=THREE; digit2<=FIVE; digit3<=FOUR; end
      16'd4536: begin digit0<=SIX; digit1<=THREE; digit2<=FIVE; digit3<=FOUR; end
      16'd4537: begin digit0<=SEVEN; digit1<=THREE; digit2<=FIVE; digit3<=FOUR; end
      16'd4538: begin digit0<=EIGHT; digit1<=THREE; digit2<=FIVE; digit3<=FOUR; end
      16'd4539: begin digit0<=NINE; digit1<=THREE; digit2<=FIVE; digit3<=FOUR; end
      16'd4540: begin digit0<=ZERO; digit1<=FOUR; digit2<=FIVE; digit3<=FOUR; end
      16'd4541: begin digit0<=ONE; digit1<=FOUR; digit2<=FIVE; digit3<=FOUR; end
      16'd4542: begin digit0<=TWO; digit1<=FOUR; digit2<=FIVE; digit3<=FOUR; end
      16'd4543: begin digit0<=THREE; digit1<=FOUR; digit2<=FIVE; digit3<=FOUR; end
      16'd4544: begin digit0<=FOUR; digit1<=FOUR; digit2<=FIVE; digit3<=FOUR; end
      16'd4545: begin digit0<=FIVE; digit1<=FOUR; digit2<=FIVE; digit3<=FOUR; end
      16'd4546: begin digit0<=SIX; digit1<=FOUR; digit2<=FIVE; digit3<=FOUR; end
      16'd4547: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FIVE; digit3<=FOUR; end
      16'd4548: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FIVE; digit3<=FOUR; end
      16'd4549: begin digit0<=NINE; digit1<=FOUR; digit2<=FIVE; digit3<=FOUR; end
      16'd4550: begin digit0<=ZERO; digit1<=FIVE; digit2<=FIVE; digit3<=FOUR; end
      16'd4551: begin digit0<=ONE; digit1<=FIVE; digit2<=FIVE; digit3<=FOUR; end
      16'd4552: begin digit0<=TWO; digit1<=FIVE; digit2<=FIVE; digit3<=FOUR; end
      16'd4553: begin digit0<=THREE; digit1<=FIVE; digit2<=FIVE; digit3<=FOUR; end
      16'd4554: begin digit0<=FOUR; digit1<=FIVE; digit2<=FIVE; digit3<=FOUR; end
      16'd4555: begin digit0<=FIVE; digit1<=FIVE; digit2<=FIVE; digit3<=FOUR; end
      16'd4556: begin digit0<=SIX; digit1<=FIVE; digit2<=FIVE; digit3<=FOUR; end
      16'd4557: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FIVE; digit3<=FOUR; end
      16'd4558: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FIVE; digit3<=FOUR; end
      16'd4559: begin digit0<=NINE; digit1<=FIVE; digit2<=FIVE; digit3<=FOUR; end
      16'd4560: begin digit0<=ZERO; digit1<=SIX; digit2<=FIVE; digit3<=FOUR; end
      16'd4561: begin digit0<=ONE; digit1<=SIX; digit2<=FIVE; digit3<=FOUR; end
      16'd4562: begin digit0<=TWO; digit1<=SIX; digit2<=FIVE; digit3<=FOUR; end
      16'd4563: begin digit0<=THREE; digit1<=SIX; digit2<=FIVE; digit3<=FOUR; end
      16'd4564: begin digit0<=FOUR; digit1<=SIX; digit2<=FIVE; digit3<=FOUR; end
      16'd4565: begin digit0<=FIVE; digit1<=SIX; digit2<=FIVE; digit3<=FOUR; end
      16'd4566: begin digit0<=SIX; digit1<=SIX; digit2<=FIVE; digit3<=FOUR; end
      16'd4567: begin digit0<=SEVEN; digit1<=SIX; digit2<=FIVE; digit3<=FOUR; end
      16'd4568: begin digit0<=EIGHT; digit1<=SIX; digit2<=FIVE; digit3<=FOUR; end
      16'd4569: begin digit0<=NINE; digit1<=SIX; digit2<=FIVE; digit3<=FOUR; end
      16'd4570: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FIVE; digit3<=FOUR; end
      16'd4571: begin digit0<=ONE; digit1<=SEVEN; digit2<=FIVE; digit3<=FOUR; end
      16'd4572: begin digit0<=TWO; digit1<=SEVEN; digit2<=FIVE; digit3<=FOUR; end
      16'd4573: begin digit0<=THREE; digit1<=SEVEN; digit2<=FIVE; digit3<=FOUR; end
      16'd4574: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FIVE; digit3<=FOUR; end
      16'd4575: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FIVE; digit3<=FOUR; end
      16'd4576: begin digit0<=SIX; digit1<=SEVEN; digit2<=FIVE; digit3<=FOUR; end
      16'd4577: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FIVE; digit3<=FOUR; end
      16'd4578: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FIVE; digit3<=FOUR; end
      16'd4579: begin digit0<=NINE; digit1<=SEVEN; digit2<=FIVE; digit3<=FOUR; end
      16'd4580: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=FOUR; end
      16'd4581: begin digit0<=ONE; digit1<=EIGHT; digit2<=FIVE; digit3<=FOUR; end
      16'd4582: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=FOUR; end
      16'd4583: begin digit0<=THREE; digit1<=EIGHT; digit2<=FIVE; digit3<=FOUR; end
      16'd4584: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FIVE; digit3<=FOUR; end
      16'd4585: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FIVE; digit3<=FOUR; end
      16'd4586: begin digit0<=SIX; digit1<=EIGHT; digit2<=FIVE; digit3<=FOUR; end
      16'd4587: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FIVE; digit3<=FOUR; end
      16'd4588: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FIVE; digit3<=FOUR; end
      16'd4589: begin digit0<=NINE; digit1<=EIGHT; digit2<=FIVE; digit3<=FOUR; end
      16'd4590: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=FOUR; end
      16'd4591: begin digit0<=ONE; digit1<=NINE; digit2<=FIVE; digit3<=FOUR; end
      16'd4592: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=FOUR; end
      16'd4593: begin digit0<=THREE; digit1<=NINE; digit2<=FIVE; digit3<=FOUR; end
      16'd4594: begin digit0<=FOUR; digit1<=NINE; digit2<=FIVE; digit3<=FOUR; end
      16'd4595: begin digit0<=FIVE; digit1<=NINE; digit2<=FIVE; digit3<=FOUR; end
      16'd4596: begin digit0<=SIX; digit1<=NINE; digit2<=FIVE; digit3<=FOUR; end
      16'd4597: begin digit0<=SEVEN; digit1<=NINE; digit2<=FIVE; digit3<=FOUR; end
      16'd4598: begin digit0<=EIGHT; digit1<=NINE; digit2<=FIVE; digit3<=FOUR; end
      16'd4599: begin digit0<=NINE; digit1<=NINE; digit2<=FIVE; digit3<=FOUR; end
	  16'd4600: begin digit0<=ZERO; digit1<=ZERO; digit2<=SIX; digit3<=FOUR; end
      16'd4601: begin digit0<=ONE; digit1<=ZERO; digit2<=SIX; digit3<=FOUR; end
      16'd4602: begin digit0<=TWO; digit1<=ZERO; digit2<=SIX; digit3<=FOUR; end
      16'd4603: begin digit0<=THREE; digit1<=ZERO; digit2<=SIX; digit3<=FOUR; end
      16'd4604: begin digit0<=FOUR; digit1<=ZERO; digit2<=SIX; digit3<=FOUR; end
      16'd4605: begin digit0<=FIVE; digit1<=ZERO; digit2<=SIX; digit3<=FOUR; end
      16'd4606: begin digit0<=SIX; digit1<=ZERO; digit2<=SIX; digit3<=FOUR; end
      16'd4607: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SIX; digit3<=FOUR; end
      16'd4608: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SIX; digit3<=FOUR; end
      16'd4609: begin digit0<=NINE; digit1<=ZERO; digit2<=SIX; digit3<=FOUR; end
      16'd4610: begin digit0<=ZERO; digit1<=ONE; digit2<=SIX; digit3<=FOUR; end
      16'd4611: begin digit0<=ONE; digit1<=ONE; digit2<=SIX; digit3<=FOUR; end
      16'd4612: begin digit0<=TWO; digit1<=ONE; digit2<=SIX; digit3<=FOUR; end
      16'd4613: begin digit0<=THREE; digit1<=ONE; digit2<=SIX; digit3<=FOUR; end
      16'd4614: begin digit0<=FOUR; digit1<=ONE; digit2<=SIX; digit3<=FOUR; end
      16'd4615: begin digit0<=FIVE; digit1<=ONE; digit2<=SIX; digit3<=FOUR; end
      16'd4616: begin digit0<=SIX; digit1<=ONE; digit2<=SIX; digit3<=FOUR; end
      16'd4617: begin digit0<=SEVEN; digit1<=ONE; digit2<=SIX; digit3<=FOUR; end
      16'd4618: begin digit0<=EIGHT; digit1<=ONE; digit2<=SIX; digit3<=FOUR; end
      16'd4619: begin digit0<=NINE; digit1<=ONE; digit2<=SIX; digit3<=FOUR; end
      16'd4620: begin digit0<=ZERO; digit1<=TWO; digit2<=SIX; digit3<=FOUR; end
      16'd4621: begin digit0<=ONE; digit1<=TWO; digit2<=SIX; digit3<=FOUR; end
      16'd4622: begin digit0<=TWO; digit1<=TWO; digit2<=SIX; digit3<=FOUR; end
      16'd4623: begin digit0<=THREE; digit1<=TWO; digit2<=SIX; digit3<=FOUR; end
      16'd4624: begin digit0<=FOUR; digit1<=TWO; digit2<=SIX; digit3<=FOUR; end
      16'd4625: begin digit0<=FIVE; digit1<=TWO; digit2<=SIX; digit3<=FOUR; end
      16'd4626: begin digit0<=SIX; digit1<=TWO; digit2<=SIX; digit3<=FOUR; end
      16'd4627: begin digit0<=SEVEN; digit1<=TWO; digit2<=SIX; digit3<=FOUR; end
      16'd4628: begin digit0<=EIGHT; digit1<=TWO; digit2<=SIX; digit3<=FOUR; end
      16'd4629: begin digit0<=NINE; digit1<=TWO; digit2<=SIX; digit3<=FOUR; end
      16'd4630: begin digit0<=ZERO; digit1<=THREE; digit2<=SIX; digit3<=FOUR; end
      16'd4631: begin digit0<=ONE; digit1<=THREE; digit2<=SIX; digit3<=FOUR; end
      16'd4632: begin digit0<=TWO; digit1<=THREE; digit2<=SIX; digit3<=FOUR; end
      16'd4633: begin digit0<=THREE; digit1<=THREE; digit2<=SIX; digit3<=FOUR; end
      16'd4634: begin digit0<=FOUR; digit1<=THREE; digit2<=SIX; digit3<=FOUR; end
      16'd4635: begin digit0<=FIVE; digit1<=THREE; digit2<=SIX; digit3<=FOUR; end
      16'd4636: begin digit0<=SIX; digit1<=THREE; digit2<=SIX; digit3<=FOUR; end
      16'd4637: begin digit0<=SEVEN; digit1<=THREE; digit2<=SIX; digit3<=FOUR; end
      16'd4638: begin digit0<=EIGHT; digit1<=THREE; digit2<=SIX; digit3<=FOUR; end
      16'd4639: begin digit0<=NINE; digit1<=THREE; digit2<=SIX; digit3<=FOUR; end
      16'd4640: begin digit0<=ZERO; digit1<=FOUR; digit2<=SIX; digit3<=FOUR; end
      16'd4641: begin digit0<=ONE; digit1<=FOUR; digit2<=SIX; digit3<=FOUR; end
      16'd4642: begin digit0<=TWO; digit1<=FOUR; digit2<=SIX; digit3<=FOUR; end
      16'd4643: begin digit0<=THREE; digit1<=FOUR; digit2<=SIX; digit3<=FOUR; end
      16'd4644: begin digit0<=FOUR; digit1<=FOUR; digit2<=SIX; digit3<=FOUR; end
      16'd4645: begin digit0<=FIVE; digit1<=FOUR; digit2<=SIX; digit3<=FOUR; end
      16'd4646: begin digit0<=SIX; digit1<=FOUR; digit2<=SIX; digit3<=FOUR; end
      16'd4647: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SIX; digit3<=FOUR; end
      16'd4648: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SIX; digit3<=FOUR; end
      16'd4649: begin digit0<=NINE; digit1<=FOUR; digit2<=SIX; digit3<=FOUR; end
      16'd4650: begin digit0<=ZERO; digit1<=FIVE; digit2<=SIX; digit3<=FOUR; end
      16'd4651: begin digit0<=ONE; digit1<=FIVE; digit2<=SIX; digit3<=FOUR; end
      16'd4652: begin digit0<=TWO; digit1<=FIVE; digit2<=SIX; digit3<=FOUR; end
      16'd4653: begin digit0<=THREE; digit1<=FIVE; digit2<=SIX; digit3<=FOUR; end
      16'd4654: begin digit0<=FOUR; digit1<=FIVE; digit2<=SIX; digit3<=FOUR; end
      16'd4655: begin digit0<=FIVE; digit1<=FIVE; digit2<=SIX; digit3<=FOUR; end
      16'd4656: begin digit0<=SIX; digit1<=FIVE; digit2<=SIX; digit3<=FOUR; end
      16'd4657: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SIX; digit3<=FOUR; end
      16'd4658: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SIX; digit3<=FOUR; end
      16'd4659: begin digit0<=NINE; digit1<=FIVE; digit2<=SIX; digit3<=FOUR; end
      16'd4660: begin digit0<=ZERO; digit1<=SIX; digit2<=SIX; digit3<=FOUR; end
      16'd4661: begin digit0<=ONE; digit1<=SIX; digit2<=SIX; digit3<=FOUR; end
      16'd4662: begin digit0<=TWO; digit1<=SIX; digit2<=SIX; digit3<=FOUR; end
      16'd4663: begin digit0<=THREE; digit1<=SIX; digit2<=SIX; digit3<=FOUR; end
      16'd4664: begin digit0<=FOUR; digit1<=SIX; digit2<=SIX; digit3<=FOUR; end
      16'd4665: begin digit0<=FIVE; digit1<=SIX; digit2<=SIX; digit3<=FOUR; end
      16'd4666: begin digit0<=SIX; digit1<=SIX; digit2<=SIX; digit3<=FOUR; end
      16'd4667: begin digit0<=SEVEN; digit1<=SIX; digit2<=SIX; digit3<=FOUR; end
      16'd4668: begin digit0<=EIGHT; digit1<=SIX; digit2<=SIX; digit3<=FOUR; end
      16'd4669: begin digit0<=NINE; digit1<=SIX; digit2<=SIX; digit3<=FOUR; end
      16'd4670: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SIX; digit3<=FOUR; end
      16'd4671: begin digit0<=ONE; digit1<=SEVEN; digit2<=SIX; digit3<=FOUR; end
      16'd4672: begin digit0<=TWO; digit1<=SEVEN; digit2<=SIX; digit3<=FOUR; end
      16'd4673: begin digit0<=THREE; digit1<=SEVEN; digit2<=SIX; digit3<=FOUR; end
      16'd4674: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SIX; digit3<=FOUR; end
      16'd4675: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SIX; digit3<=FOUR; end
      16'd4676: begin digit0<=SIX; digit1<=SEVEN; digit2<=SIX; digit3<=FOUR; end
      16'd4677: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SIX; digit3<=FOUR; end
      16'd4678: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SIX; digit3<=FOUR; end
      16'd4679: begin digit0<=NINE; digit1<=SEVEN; digit2<=SIX; digit3<=FOUR; end
      16'd4680: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=FOUR; end
      16'd4681: begin digit0<=ONE; digit1<=EIGHT; digit2<=SIX; digit3<=FOUR; end
      16'd4682: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=FOUR; end
      16'd4683: begin digit0<=THREE; digit1<=EIGHT; digit2<=SIX; digit3<=FOUR; end
      16'd4684: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SIX; digit3<=FOUR; end
      16'd4685: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SIX; digit3<=FOUR; end
      16'd4686: begin digit0<=SIX; digit1<=EIGHT; digit2<=SIX; digit3<=FOUR; end
      16'd4687: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SIX; digit3<=FOUR; end
      16'd4688: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SIX; digit3<=FOUR; end
      16'd4689: begin digit0<=NINE; digit1<=EIGHT; digit2<=SIX; digit3<=FOUR; end
      16'd4690: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=FOUR; end
      16'd4691: begin digit0<=ONE; digit1<=NINE; digit2<=SIX; digit3<=FOUR; end
      16'd4692: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=FOUR; end
      16'd4693: begin digit0<=THREE; digit1<=NINE; digit2<=SIX; digit3<=FOUR; end
      16'd4694: begin digit0<=FOUR; digit1<=NINE; digit2<=SIX; digit3<=FOUR; end
      16'd4695: begin digit0<=FIVE; digit1<=NINE; digit2<=SIX; digit3<=FOUR; end
      16'd4696: begin digit0<=SIX; digit1<=NINE; digit2<=SIX; digit3<=FOUR; end
      16'd4697: begin digit0<=SEVEN; digit1<=NINE; digit2<=SIX; digit3<=FOUR; end
      16'd4698: begin digit0<=EIGHT; digit1<=NINE; digit2<=SIX; digit3<=FOUR; end
      16'd4699: begin digit0<=NINE; digit1<=NINE; digit2<=SIX; digit3<=FOUR; end
	  16'd4700: begin digit0<=ZERO; digit1<=ZERO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4701: begin digit0<=ONE; digit1<=ZERO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4702: begin digit0<=TWO; digit1<=ZERO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4703: begin digit0<=THREE; digit1<=ZERO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4704: begin digit0<=FOUR; digit1<=ZERO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4705: begin digit0<=FIVE; digit1<=ZERO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4706: begin digit0<=SIX; digit1<=ZERO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4707: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4708: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4709: begin digit0<=NINE; digit1<=ZERO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4710: begin digit0<=ZERO; digit1<=ONE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4711: begin digit0<=ONE; digit1<=ONE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4712: begin digit0<=TWO; digit1<=ONE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4713: begin digit0<=THREE; digit1<=ONE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4714: begin digit0<=FOUR; digit1<=ONE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4715: begin digit0<=FIVE; digit1<=ONE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4716: begin digit0<=SIX; digit1<=ONE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4717: begin digit0<=SEVEN; digit1<=ONE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4718: begin digit0<=EIGHT; digit1<=ONE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4719: begin digit0<=NINE; digit1<=ONE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4720: begin digit0<=ZERO; digit1<=TWO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4721: begin digit0<=ONE; digit1<=TWO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4722: begin digit0<=TWO; digit1<=TWO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4723: begin digit0<=THREE; digit1<=TWO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4724: begin digit0<=FOUR; digit1<=TWO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4725: begin digit0<=FIVE; digit1<=TWO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4726: begin digit0<=SIX; digit1<=TWO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4727: begin digit0<=SEVEN; digit1<=TWO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4728: begin digit0<=EIGHT; digit1<=TWO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4729: begin digit0<=NINE; digit1<=TWO; digit2<=SEVEN; digit3<=FOUR; end
      16'd4730: begin digit0<=ZERO; digit1<=THREE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4731: begin digit0<=ONE; digit1<=THREE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4732: begin digit0<=TWO; digit1<=THREE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4733: begin digit0<=THREE; digit1<=THREE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4734: begin digit0<=FOUR; digit1<=THREE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4735: begin digit0<=FIVE; digit1<=THREE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4736: begin digit0<=SIX; digit1<=THREE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4737: begin digit0<=SEVEN; digit1<=THREE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4738: begin digit0<=EIGHT; digit1<=THREE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4739: begin digit0<=NINE; digit1<=THREE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4740: begin digit0<=ZERO; digit1<=FOUR; digit2<=SEVEN; digit3<=FOUR; end
      16'd4741: begin digit0<=ONE; digit1<=FOUR; digit2<=SEVEN; digit3<=FOUR; end
      16'd4742: begin digit0<=TWO; digit1<=FOUR; digit2<=SEVEN; digit3<=FOUR; end
      16'd4743: begin digit0<=THREE; digit1<=FOUR; digit2<=SEVEN; digit3<=FOUR; end
      16'd4744: begin digit0<=FOUR; digit1<=FOUR; digit2<=SEVEN; digit3<=FOUR; end
      16'd4745: begin digit0<=FIVE; digit1<=FOUR; digit2<=SEVEN; digit3<=FOUR; end
      16'd4746: begin digit0<=SIX; digit1<=FOUR; digit2<=SEVEN; digit3<=FOUR; end
      16'd4747: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SEVEN; digit3<=FOUR; end
      16'd4748: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SEVEN; digit3<=FOUR; end
      16'd4749: begin digit0<=NINE; digit1<=FOUR; digit2<=SEVEN; digit3<=FOUR; end
      16'd4750: begin digit0<=ZERO; digit1<=FIVE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4751: begin digit0<=ONE; digit1<=FIVE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4752: begin digit0<=TWO; digit1<=FIVE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4753: begin digit0<=THREE; digit1<=FIVE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4754: begin digit0<=FOUR; digit1<=FIVE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4755: begin digit0<=FIVE; digit1<=FIVE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4756: begin digit0<=SIX; digit1<=FIVE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4757: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4758: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4759: begin digit0<=NINE; digit1<=FIVE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4760: begin digit0<=ZERO; digit1<=SIX; digit2<=SEVEN; digit3<=FOUR; end
      16'd4761: begin digit0<=ONE; digit1<=SIX; digit2<=SEVEN; digit3<=FOUR; end
      16'd4762: begin digit0<=TWO; digit1<=SIX; digit2<=SEVEN; digit3<=FOUR; end
      16'd4763: begin digit0<=THREE; digit1<=SIX; digit2<=SEVEN; digit3<=FOUR; end
      16'd4764: begin digit0<=FOUR; digit1<=SIX; digit2<=SEVEN; digit3<=FOUR; end
      16'd4765: begin digit0<=FIVE; digit1<=SIX; digit2<=SEVEN; digit3<=FOUR; end
      16'd4766: begin digit0<=SIX; digit1<=SIX; digit2<=SEVEN; digit3<=FOUR; end
      16'd4767: begin digit0<=SEVEN; digit1<=SIX; digit2<=SEVEN; digit3<=FOUR; end
      16'd4768: begin digit0<=EIGHT; digit1<=SIX; digit2<=SEVEN; digit3<=FOUR; end
      16'd4769: begin digit0<=NINE; digit1<=SIX; digit2<=SEVEN; digit3<=FOUR; end
      16'd4770: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SEVEN; digit3<=FOUR; end
      16'd4771: begin digit0<=ONE; digit1<=SEVEN; digit2<=SEVEN; digit3<=FOUR; end
      16'd4772: begin digit0<=TWO; digit1<=SEVEN; digit2<=SEVEN; digit3<=FOUR; end
      16'd4773: begin digit0<=THREE; digit1<=SEVEN; digit2<=SEVEN; digit3<=FOUR; end
      16'd4774: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SEVEN; digit3<=FOUR; end
      16'd4775: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SEVEN; digit3<=FOUR; end
      16'd4776: begin digit0<=SIX; digit1<=SEVEN; digit2<=SEVEN; digit3<=FOUR; end
      16'd4777: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SEVEN; digit3<=FOUR; end
      16'd4778: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SEVEN; digit3<=FOUR; end
      16'd4779: begin digit0<=NINE; digit1<=SEVEN; digit2<=SEVEN; digit3<=FOUR; end
      16'd4780: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=FOUR; end
      16'd4781: begin digit0<=ONE; digit1<=EIGHT; digit2<=SEVEN; digit3<=FOUR; end
      16'd4782: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=FOUR; end
      16'd4783: begin digit0<=THREE; digit1<=EIGHT; digit2<=SEVEN; digit3<=FOUR; end
      16'd4784: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SEVEN; digit3<=FOUR; end
      16'd4785: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SEVEN; digit3<=FOUR; end
      16'd4786: begin digit0<=SIX; digit1<=EIGHT; digit2<=SEVEN; digit3<=FOUR; end
      16'd4787: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SEVEN; digit3<=FOUR; end
      16'd4788: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SEVEN; digit3<=FOUR; end
      16'd4789: begin digit0<=NINE; digit1<=EIGHT; digit2<=SEVEN; digit3<=FOUR; end
      16'd4790: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4791: begin digit0<=ONE; digit1<=NINE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4792: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4793: begin digit0<=THREE; digit1<=NINE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4794: begin digit0<=FOUR; digit1<=NINE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4795: begin digit0<=FIVE; digit1<=NINE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4796: begin digit0<=SIX; digit1<=NINE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4797: begin digit0<=SEVEN; digit1<=NINE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4798: begin digit0<=EIGHT; digit1<=NINE; digit2<=SEVEN; digit3<=FOUR; end
      16'd4799: begin digit0<=NINE; digit1<=NINE; digit2<=SEVEN; digit3<=FOUR; end
	  16'd4800: begin digit0<=ZERO; digit1<=ZERO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4801: begin digit0<=ONE; digit1<=ZERO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4802: begin digit0<=TWO; digit1<=ZERO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4803: begin digit0<=THREE; digit1<=ZERO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4804: begin digit0<=FOUR; digit1<=ZERO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4805: begin digit0<=FIVE; digit1<=ZERO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4806: begin digit0<=SIX; digit1<=ZERO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4807: begin digit0<=SEVEN; digit1<=ZERO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4808: begin digit0<=EIGHT; digit1<=ZERO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4809: begin digit0<=NINE; digit1<=ZERO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4810: begin digit0<=ZERO; digit1<=ONE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4811: begin digit0<=ONE; digit1<=ONE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4812: begin digit0<=TWO; digit1<=ONE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4813: begin digit0<=THREE; digit1<=ONE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4814: begin digit0<=FOUR; digit1<=ONE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4815: begin digit0<=FIVE; digit1<=ONE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4816: begin digit0<=SIX; digit1<=ONE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4817: begin digit0<=SEVEN; digit1<=ONE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4818: begin digit0<=EIGHT; digit1<=ONE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4819: begin digit0<=NINE; digit1<=ONE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4820: begin digit0<=ZERO; digit1<=TWO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4821: begin digit0<=ONE; digit1<=TWO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4822: begin digit0<=TWO; digit1<=TWO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4823: begin digit0<=THREE; digit1<=TWO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4824: begin digit0<=FOUR; digit1<=TWO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4825: begin digit0<=FIVE; digit1<=TWO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4826: begin digit0<=SIX; digit1<=TWO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4827: begin digit0<=SEVEN; digit1<=TWO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4828: begin digit0<=EIGHT; digit1<=TWO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4829: begin digit0<=NINE; digit1<=TWO; digit2<=EIGHT; digit3<=FOUR; end
      16'd4830: begin digit0<=ZERO; digit1<=THREE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4831: begin digit0<=ONE; digit1<=THREE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4832: begin digit0<=TWO; digit1<=THREE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4833: begin digit0<=THREE; digit1<=THREE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4834: begin digit0<=FOUR; digit1<=THREE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4835: begin digit0<=FIVE; digit1<=THREE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4836: begin digit0<=SIX; digit1<=THREE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4837: begin digit0<=SEVEN; digit1<=THREE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4838: begin digit0<=EIGHT; digit1<=THREE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4839: begin digit0<=NINE; digit1<=THREE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4840: begin digit0<=ZERO; digit1<=FOUR; digit2<=EIGHT; digit3<=FOUR; end
      16'd4841: begin digit0<=ONE; digit1<=FOUR; digit2<=EIGHT; digit3<=FOUR; end
      16'd4842: begin digit0<=TWO; digit1<=FOUR; digit2<=EIGHT; digit3<=FOUR; end
      16'd4843: begin digit0<=THREE; digit1<=FOUR; digit2<=EIGHT; digit3<=FOUR; end
      16'd4844: begin digit0<=FOUR; digit1<=FOUR; digit2<=EIGHT; digit3<=FOUR; end
      16'd4845: begin digit0<=FIVE; digit1<=FOUR; digit2<=EIGHT; digit3<=FOUR; end
      16'd4846: begin digit0<=SIX; digit1<=FOUR; digit2<=EIGHT; digit3<=FOUR; end
      16'd4847: begin digit0<=SEVEN; digit1<=FOUR; digit2<=EIGHT; digit3<=FOUR; end
      16'd4848: begin digit0<=EIGHT; digit1<=FOUR; digit2<=EIGHT; digit3<=FOUR; end
      16'd4849: begin digit0<=NINE; digit1<=FOUR; digit2<=EIGHT; digit3<=FOUR; end
      16'd4850: begin digit0<=ZERO; digit1<=FIVE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4851: begin digit0<=ONE; digit1<=FIVE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4852: begin digit0<=TWO; digit1<=FIVE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4853: begin digit0<=THREE; digit1<=FIVE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4854: begin digit0<=FOUR; digit1<=FIVE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4855: begin digit0<=FIVE; digit1<=FIVE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4856: begin digit0<=SIX; digit1<=FIVE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4857: begin digit0<=SEVEN; digit1<=FIVE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4858: begin digit0<=EIGHT; digit1<=FIVE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4859: begin digit0<=NINE; digit1<=FIVE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4860: begin digit0<=ZERO; digit1<=SIX; digit2<=EIGHT; digit3<=FOUR; end
      16'd4861: begin digit0<=ONE; digit1<=SIX; digit2<=EIGHT; digit3<=FOUR; end
      16'd4862: begin digit0<=TWO; digit1<=SIX; digit2<=EIGHT; digit3<=FOUR; end
      16'd4863: begin digit0<=THREE; digit1<=SIX; digit2<=EIGHT; digit3<=FOUR; end
      16'd4864: begin digit0<=FOUR; digit1<=SIX; digit2<=EIGHT; digit3<=FOUR; end
      16'd4865: begin digit0<=FIVE; digit1<=SIX; digit2<=EIGHT; digit3<=FOUR; end
      16'd4866: begin digit0<=SIX; digit1<=SIX; digit2<=EIGHT; digit3<=FOUR; end
      16'd4867: begin digit0<=SEVEN; digit1<=SIX; digit2<=EIGHT; digit3<=FOUR; end
      16'd4868: begin digit0<=EIGHT; digit1<=SIX; digit2<=EIGHT; digit3<=FOUR; end
      16'd4869: begin digit0<=NINE; digit1<=SIX; digit2<=EIGHT; digit3<=FOUR; end
      16'd4870: begin digit0<=ZERO; digit1<=SEVEN; digit2<=EIGHT; digit3<=FOUR; end
      16'd4871: begin digit0<=ONE; digit1<=SEVEN; digit2<=EIGHT; digit3<=FOUR; end
      16'd4872: begin digit0<=TWO; digit1<=SEVEN; digit2<=EIGHT; digit3<=FOUR; end
      16'd4873: begin digit0<=THREE; digit1<=SEVEN; digit2<=EIGHT; digit3<=FOUR; end
      16'd4874: begin digit0<=FOUR; digit1<=SEVEN; digit2<=EIGHT; digit3<=FOUR; end
      16'd4875: begin digit0<=FIVE; digit1<=SEVEN; digit2<=EIGHT; digit3<=FOUR; end
      16'd4876: begin digit0<=SIX; digit1<=SEVEN; digit2<=EIGHT; digit3<=FOUR; end
      16'd4877: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=EIGHT; digit3<=FOUR; end
      16'd4878: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=EIGHT; digit3<=FOUR; end
      16'd4879: begin digit0<=NINE; digit1<=SEVEN; digit2<=EIGHT; digit3<=FOUR; end
      16'd4880: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=FOUR; end
      16'd4881: begin digit0<=ONE; digit1<=EIGHT; digit2<=EIGHT; digit3<=FOUR; end
      16'd4882: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=FOUR; end
      16'd4883: begin digit0<=THREE; digit1<=EIGHT; digit2<=EIGHT; digit3<=FOUR; end
      16'd4884: begin digit0<=FOUR; digit1<=EIGHT; digit2<=EIGHT; digit3<=FOUR; end
      16'd4885: begin digit0<=FIVE; digit1<=EIGHT; digit2<=EIGHT; digit3<=FOUR; end
      16'd4886: begin digit0<=SIX; digit1<=EIGHT; digit2<=EIGHT; digit3<=FOUR; end
      16'd4887: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=EIGHT; digit3<=FOUR; end
      16'd4888: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=EIGHT; digit3<=FOUR; end
      16'd4889: begin digit0<=NINE; digit1<=EIGHT; digit2<=EIGHT; digit3<=FOUR; end
      16'd4890: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4891: begin digit0<=ONE; digit1<=NINE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4892: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4893: begin digit0<=THREE; digit1<=NINE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4894: begin digit0<=FOUR; digit1<=NINE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4895: begin digit0<=FIVE; digit1<=NINE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4896: begin digit0<=SIX; digit1<=NINE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4897: begin digit0<=SEVEN; digit1<=NINE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4898: begin digit0<=EIGHT; digit1<=NINE; digit2<=EIGHT; digit3<=FOUR; end
      16'd4899: begin digit0<=NINE; digit1<=NINE; digit2<=EIGHT; digit3<=FOUR; end
	  16'd4900: begin digit0<=ZERO; digit1<=ZERO; digit2<=NINE; digit3<=FOUR; end
      16'd4901: begin digit0<=ONE; digit1<=ZERO; digit2<=NINE; digit3<=FOUR; end
      16'd4902: begin digit0<=TWO; digit1<=ZERO; digit2<=NINE; digit3<=FOUR; end
      16'd4903: begin digit0<=THREE; digit1<=ZERO; digit2<=NINE; digit3<=FOUR; end
      16'd4904: begin digit0<=FOUR; digit1<=ZERO; digit2<=NINE; digit3<=FOUR; end
      16'd4905: begin digit0<=FIVE; digit1<=ZERO; digit2<=NINE; digit3<=FOUR; end
      16'd4906: begin digit0<=SIX; digit1<=ZERO; digit2<=NINE; digit3<=FOUR; end
      16'd4907: begin digit0<=SEVEN; digit1<=ZERO; digit2<=NINE; digit3<=FOUR; end
      16'd4908: begin digit0<=EIGHT; digit1<=ZERO; digit2<=NINE; digit3<=FOUR; end
      16'd4909: begin digit0<=NINE; digit1<=ZERO; digit2<=NINE; digit3<=FOUR; end
      16'd4910: begin digit0<=ZERO; digit1<=ONE; digit2<=NINE; digit3<=FOUR; end
      16'd4911: begin digit0<=ONE; digit1<=ONE; digit2<=NINE; digit3<=FOUR; end
      16'd4912: begin digit0<=TWO; digit1<=ONE; digit2<=NINE; digit3<=FOUR; end
      16'd4913: begin digit0<=THREE; digit1<=ONE; digit2<=NINE; digit3<=FOUR; end
      16'd4914: begin digit0<=FOUR; digit1<=ONE; digit2<=NINE; digit3<=FOUR; end
      16'd4915: begin digit0<=FIVE; digit1<=ONE; digit2<=NINE; digit3<=FOUR; end
      16'd4916: begin digit0<=SIX; digit1<=ONE; digit2<=NINE; digit3<=FOUR; end
      16'd4917: begin digit0<=SEVEN; digit1<=ONE; digit2<=NINE; digit3<=FOUR; end
      16'd4918: begin digit0<=EIGHT; digit1<=ONE; digit2<=NINE; digit3<=FOUR; end
      16'd4919: begin digit0<=NINE; digit1<=ONE; digit2<=NINE; digit3<=FOUR; end
      16'd4920: begin digit0<=ZERO; digit1<=TWO; digit2<=NINE; digit3<=FOUR; end
      16'd4921: begin digit0<=ONE; digit1<=TWO; digit2<=NINE; digit3<=FOUR; end
      16'd4922: begin digit0<=TWO; digit1<=TWO; digit2<=NINE; digit3<=FOUR; end
      16'd4923: begin digit0<=THREE; digit1<=TWO; digit2<=NINE; digit3<=FOUR; end
      16'd4924: begin digit0<=FOUR; digit1<=TWO; digit2<=NINE; digit3<=FOUR; end
      16'd4925: begin digit0<=FIVE; digit1<=TWO; digit2<=NINE; digit3<=FOUR; end
      16'd4926: begin digit0<=SIX; digit1<=TWO; digit2<=NINE; digit3<=FOUR; end
      16'd4927: begin digit0<=SEVEN; digit1<=TWO; digit2<=NINE; digit3<=FOUR; end
      16'd4928: begin digit0<=EIGHT; digit1<=TWO; digit2<=NINE; digit3<=FOUR; end
      16'd4929: begin digit0<=NINE; digit1<=TWO; digit2<=NINE; digit3<=FOUR; end
      16'd4930: begin digit0<=ZERO; digit1<=THREE; digit2<=NINE; digit3<=FOUR; end
      16'd4931: begin digit0<=ONE; digit1<=THREE; digit2<=NINE; digit3<=FOUR; end
      16'd4932: begin digit0<=TWO; digit1<=THREE; digit2<=NINE; digit3<=FOUR; end
      16'd4933: begin digit0<=THREE; digit1<=THREE; digit2<=NINE; digit3<=FOUR; end
      16'd4934: begin digit0<=FOUR; digit1<=THREE; digit2<=NINE; digit3<=FOUR; end
      16'd4935: begin digit0<=FIVE; digit1<=THREE; digit2<=NINE; digit3<=FOUR; end
      16'd4936: begin digit0<=SIX; digit1<=THREE; digit2<=NINE; digit3<=FOUR; end
      16'd4937: begin digit0<=SEVEN; digit1<=THREE; digit2<=NINE; digit3<=FOUR; end
      16'd4938: begin digit0<=EIGHT; digit1<=THREE; digit2<=NINE; digit3<=FOUR; end
      16'd4939: begin digit0<=NINE; digit1<=THREE; digit2<=NINE; digit3<=FOUR; end
      16'd4940: begin digit0<=ZERO; digit1<=FOUR; digit2<=NINE; digit3<=FOUR; end
      16'd4941: begin digit0<=ONE; digit1<=FOUR; digit2<=NINE; digit3<=FOUR; end
      16'd4942: begin digit0<=TWO; digit1<=FOUR; digit2<=NINE; digit3<=FOUR; end
      16'd4943: begin digit0<=THREE; digit1<=FOUR; digit2<=NINE; digit3<=FOUR; end
      16'd4944: begin digit0<=FOUR; digit1<=FOUR; digit2<=NINE; digit3<=FOUR; end
      16'd4945: begin digit0<=FIVE; digit1<=FOUR; digit2<=NINE; digit3<=FOUR; end
      16'd4946: begin digit0<=SIX; digit1<=FOUR; digit2<=NINE; digit3<=FOUR; end
      16'd4947: begin digit0<=SEVEN; digit1<=FOUR; digit2<=NINE; digit3<=FOUR; end
      16'd4948: begin digit0<=EIGHT; digit1<=FOUR; digit2<=NINE; digit3<=FOUR; end
      16'd4949: begin digit0<=NINE; digit1<=FOUR; digit2<=NINE; digit3<=FOUR; end
      16'd4950: begin digit0<=ZERO; digit1<=FIVE; digit2<=NINE; digit3<=FOUR; end
      16'd4951: begin digit0<=ONE; digit1<=FIVE; digit2<=NINE; digit3<=FOUR; end
      16'd4952: begin digit0<=TWO; digit1<=FIVE; digit2<=NINE; digit3<=FOUR; end
      16'd4953: begin digit0<=THREE; digit1<=FIVE; digit2<=NINE; digit3<=FOUR; end
      16'd4954: begin digit0<=FOUR; digit1<=FIVE; digit2<=NINE; digit3<=FOUR; end
      16'd4955: begin digit0<=FIVE; digit1<=FIVE; digit2<=NINE; digit3<=FOUR; end
      16'd4956: begin digit0<=SIX; digit1<=FIVE; digit2<=NINE; digit3<=FOUR; end
      16'd4957: begin digit0<=SEVEN; digit1<=FIVE; digit2<=NINE; digit3<=FOUR; end
      16'd4958: begin digit0<=EIGHT; digit1<=FIVE; digit2<=NINE; digit3<=FOUR; end
      16'd4959: begin digit0<=NINE; digit1<=FIVE; digit2<=NINE; digit3<=FOUR; end
      16'd4960: begin digit0<=ZERO; digit1<=SIX; digit2<=NINE; digit3<=FOUR; end
      16'd4961: begin digit0<=ONE; digit1<=SIX; digit2<=NINE; digit3<=FOUR; end
      16'd4962: begin digit0<=TWO; digit1<=SIX; digit2<=NINE; digit3<=FOUR; end
      16'd4963: begin digit0<=THREE; digit1<=SIX; digit2<=NINE; digit3<=FOUR; end
      16'd4964: begin digit0<=FOUR; digit1<=SIX; digit2<=NINE; digit3<=FOUR; end
      16'd4965: begin digit0<=FIVE; digit1<=SIX; digit2<=NINE; digit3<=FOUR; end
      16'd4966: begin digit0<=SIX; digit1<=SIX; digit2<=NINE; digit3<=FOUR; end
      16'd4967: begin digit0<=SEVEN; digit1<=SIX; digit2<=NINE; digit3<=FOUR; end
      16'd4968: begin digit0<=EIGHT; digit1<=SIX; digit2<=NINE; digit3<=FOUR; end
      16'd4969: begin digit0<=NINE; digit1<=SIX; digit2<=NINE; digit3<=FOUR; end
      16'd4970: begin digit0<=ZERO; digit1<=SEVEN; digit2<=NINE; digit3<=FOUR; end
      16'd4971: begin digit0<=ONE; digit1<=SEVEN; digit2<=NINE; digit3<=FOUR; end
      16'd4972: begin digit0<=TWO; digit1<=SEVEN; digit2<=NINE; digit3<=FOUR; end
      16'd4973: begin digit0<=THREE; digit1<=SEVEN; digit2<=NINE; digit3<=FOUR; end
      16'd4974: begin digit0<=FOUR; digit1<=SEVEN; digit2<=NINE; digit3<=FOUR; end
      16'd4975: begin digit0<=FIVE; digit1<=SEVEN; digit2<=NINE; digit3<=FOUR; end
      16'd4976: begin digit0<=SIX; digit1<=SEVEN; digit2<=NINE; digit3<=FOUR; end
      16'd4977: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=NINE; digit3<=FOUR; end
      16'd4978: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=NINE; digit3<=FOUR; end
      16'd4979: begin digit0<=NINE; digit1<=SEVEN; digit2<=NINE; digit3<=FOUR; end
      16'd4980: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=FOUR; end
      16'd4981: begin digit0<=ONE; digit1<=EIGHT; digit2<=NINE; digit3<=FOUR; end
      16'd4982: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=FOUR; end
      16'd4983: begin digit0<=THREE; digit1<=EIGHT; digit2<=NINE; digit3<=FOUR; end
      16'd4984: begin digit0<=FOUR; digit1<=EIGHT; digit2<=NINE; digit3<=FOUR; end
      16'd4985: begin digit0<=FIVE; digit1<=EIGHT; digit2<=NINE; digit3<=FOUR; end
      16'd4986: begin digit0<=SIX; digit1<=EIGHT; digit2<=NINE; digit3<=FOUR; end
      16'd4987: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=NINE; digit3<=FOUR; end
      16'd4988: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=NINE; digit3<=FOUR; end
      16'd4989: begin digit0<=NINE; digit1<=EIGHT; digit2<=NINE; digit3<=FOUR; end
      16'd4990: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=FOUR; end
      16'd4991: begin digit0<=ONE; digit1<=NINE; digit2<=NINE; digit3<=FOUR; end
      16'd4992: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=FOUR; end
      16'd4993: begin digit0<=THREE; digit1<=NINE; digit2<=NINE; digit3<=FOUR; end
      16'd4994: begin digit0<=FOUR; digit1<=NINE; digit2<=NINE; digit3<=FOUR; end
      16'd4995: begin digit0<=FIVE; digit1<=NINE; digit2<=NINE; digit3<=FOUR; end
      16'd4996: begin digit0<=SIX; digit1<=NINE; digit2<=NINE; digit3<=FOUR; end
      16'd4997: begin digit0<=SEVEN; digit1<=NINE; digit2<=NINE; digit3<=FOUR; end
      16'd4998: begin digit0<=EIGHT; digit1<=NINE; digit2<=NINE; digit3<=FOUR; end
      16'd4999: begin digit0<=NINE; digit1<=NINE; digit2<=NINE; digit3<=FOUR; end
	  16'd5000: begin digit0<=ZERO; digit1<=ZERO; digit2<=ZERO; digit3<=FIVE; end
      16'd5001: begin digit0<=ONE; digit1<=ZERO; digit2<=ZERO; digit3<=FIVE; end
      16'd5002: begin digit0<=TWO; digit1<=ZERO; digit2<=ZERO; digit3<=FIVE; end
      16'd5003: begin digit0<=THREE; digit1<=ZERO; digit2<=ZERO; digit3<=FIVE; end
      16'd5004: begin digit0<=FOUR; digit1<=ZERO; digit2<=ZERO; digit3<=FIVE; end
      16'd5005: begin digit0<=FIVE; digit1<=ZERO; digit2<=ZERO; digit3<=FIVE; end
      16'd5006: begin digit0<=SIX; digit1<=ZERO; digit2<=ZERO; digit3<=FIVE; end
      16'd5007: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ZERO; digit3<=FIVE; end
      16'd5008: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ZERO; digit3<=FIVE; end
      16'd5009: begin digit0<=NINE; digit1<=ZERO; digit2<=ZERO; digit3<=FIVE; end
      16'd5010: begin digit0<=ZERO; digit1<=ONE; digit2<=ZERO; digit3<=FIVE; end
      16'd5011: begin digit0<=ONE; digit1<=ONE; digit2<=ZERO; digit3<=FIVE; end
      16'd5012: begin digit0<=TWO; digit1<=ONE; digit2<=ZERO; digit3<=FIVE; end
      16'd5013: begin digit0<=THREE; digit1<=ONE; digit2<=ZERO; digit3<=FIVE; end
      16'd5014: begin digit0<=FOUR; digit1<=ONE; digit2<=ZERO; digit3<=FIVE; end
      16'd5015: begin digit0<=FIVE; digit1<=ONE; digit2<=ZERO; digit3<=FIVE; end
      16'd5016: begin digit0<=SIX; digit1<=ONE; digit2<=ZERO; digit3<=FIVE; end
      16'd5017: begin digit0<=SEVEN; digit1<=ONE; digit2<=ZERO; digit3<=FIVE; end
      16'd5018: begin digit0<=EIGHT; digit1<=ONE; digit2<=ZERO; digit3<=FIVE; end
      16'd5019: begin digit0<=NINE; digit1<=ONE; digit2<=ZERO; digit3<=FIVE; end
      16'd5020: begin digit0<=ZERO; digit1<=TWO; digit2<=ZERO; digit3<=FIVE; end
      16'd5021: begin digit0<=ONE; digit1<=TWO; digit2<=ZERO; digit3<=FIVE; end
      16'd5022: begin digit0<=TWO; digit1<=TWO; digit2<=ZERO; digit3<=FIVE; end
      16'd5023: begin digit0<=THREE; digit1<=TWO; digit2<=ZERO; digit3<=FIVE; end
      16'd5024: begin digit0<=FOUR; digit1<=TWO; digit2<=ZERO; digit3<=FIVE; end
      16'd5025: begin digit0<=FIVE; digit1<=TWO; digit2<=ZERO; digit3<=FIVE; end
      16'd5026: begin digit0<=SIX; digit1<=TWO; digit2<=ZERO; digit3<=FIVE; end
      16'd5027: begin digit0<=SEVEN; digit1<=TWO; digit2<=ZERO; digit3<=FIVE; end
      16'd5028: begin digit0<=EIGHT; digit1<=TWO; digit2<=ZERO; digit3<=FIVE; end
      16'd5029: begin digit0<=NINE; digit1<=TWO; digit2<=ZERO; digit3<=FIVE; end
      16'd5030: begin digit0<=ZERO; digit1<=THREE; digit2<=ZERO; digit3<=FIVE; end
      16'd5031: begin digit0<=ONE; digit1<=THREE; digit2<=ZERO; digit3<=FIVE; end
      16'd5032: begin digit0<=TWO; digit1<=THREE; digit2<=ZERO; digit3<=FIVE; end
      16'd5033: begin digit0<=THREE; digit1<=THREE; digit2<=ZERO; digit3<=FIVE; end
      16'd5034: begin digit0<=FOUR; digit1<=THREE; digit2<=ZERO; digit3<=FIVE; end
      16'd5035: begin digit0<=FIVE; digit1<=THREE; digit2<=ZERO; digit3<=FIVE; end
      16'd5036: begin digit0<=SIX; digit1<=THREE; digit2<=ZERO; digit3<=FIVE; end
      16'd5037: begin digit0<=SEVEN; digit1<=THREE; digit2<=ZERO; digit3<=FIVE; end
      16'd5038: begin digit0<=EIGHT; digit1<=THREE; digit2<=ZERO; digit3<=FIVE; end
      16'd5039: begin digit0<=NINE; digit1<=THREE; digit2<=ZERO; digit3<=FIVE; end
      16'd5040: begin digit0<=ZERO; digit1<=FOUR; digit2<=ZERO; digit3<=FIVE; end
      16'd5041: begin digit0<=ONE; digit1<=FOUR; digit2<=ZERO; digit3<=FIVE; end
      16'd5042: begin digit0<=TWO; digit1<=FOUR; digit2<=ZERO; digit3<=FIVE; end
      16'd5043: begin digit0<=THREE; digit1<=FOUR; digit2<=ZERO; digit3<=FIVE; end
      16'd5044: begin digit0<=FOUR; digit1<=FOUR; digit2<=ZERO; digit3<=FIVE; end
      16'd5045: begin digit0<=FIVE; digit1<=FOUR; digit2<=ZERO; digit3<=FIVE; end
      16'd5046: begin digit0<=SIX; digit1<=FOUR; digit2<=ZERO; digit3<=FIVE; end
      16'd5047: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ZERO; digit3<=FIVE; end
      16'd5048: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ZERO; digit3<=FIVE; end
      16'd5049: begin digit0<=NINE; digit1<=FOUR; digit2<=ZERO; digit3<=FIVE; end
      16'd5050: begin digit0<=ZERO; digit1<=FIVE; digit2<=ZERO; digit3<=FIVE; end
      16'd5051: begin digit0<=ONE; digit1<=FIVE; digit2<=ZERO; digit3<=FIVE; end
      16'd5052: begin digit0<=TWO; digit1<=FIVE; digit2<=ZERO; digit3<=FIVE; end
      16'd5053: begin digit0<=THREE; digit1<=FIVE; digit2<=ZERO; digit3<=FIVE; end
      16'd5054: begin digit0<=FOUR; digit1<=FIVE; digit2<=ZERO; digit3<=FIVE; end
      16'd5055: begin digit0<=FIVE; digit1<=FIVE; digit2<=ZERO; digit3<=FIVE; end
      16'd5056: begin digit0<=SIX; digit1<=FIVE; digit2<=ZERO; digit3<=FIVE; end
      16'd5057: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ZERO; digit3<=FIVE; end
      16'd5058: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ZERO; digit3<=FIVE; end
      16'd5059: begin digit0<=NINE; digit1<=FIVE; digit2<=ZERO; digit3<=FIVE; end
      16'd5060: begin digit0<=ZERO; digit1<=SIX; digit2<=ZERO; digit3<=FIVE; end
      16'd5061: begin digit0<=ONE; digit1<=SIX; digit2<=ZERO; digit3<=FIVE; end
      16'd5062: begin digit0<=TWO; digit1<=SIX; digit2<=ZERO; digit3<=FIVE; end
      16'd5063: begin digit0<=THREE; digit1<=SIX; digit2<=ZERO; digit3<=FIVE; end
      16'd5064: begin digit0<=FOUR; digit1<=SIX; digit2<=ZERO; digit3<=FIVE; end
      16'd5065: begin digit0<=FIVE; digit1<=SIX; digit2<=ZERO; digit3<=FIVE; end
      16'd5066: begin digit0<=SIX; digit1<=SIX; digit2<=ZERO; digit3<=FIVE; end
      16'd5067: begin digit0<=SEVEN; digit1<=SIX; digit2<=ZERO; digit3<=FIVE; end
      16'd5068: begin digit0<=EIGHT; digit1<=SIX; digit2<=ZERO; digit3<=FIVE; end
      16'd5069: begin digit0<=NINE; digit1<=SIX; digit2<=ZERO; digit3<=FIVE; end
      16'd5070: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ZERO; digit3<=FIVE; end
      16'd5071: begin digit0<=ONE; digit1<=SEVEN; digit2<=ZERO; digit3<=FIVE; end
      16'd5072: begin digit0<=TWO; digit1<=SEVEN; digit2<=ZERO; digit3<=FIVE; end
      16'd5073: begin digit0<=THREE; digit1<=SEVEN; digit2<=ZERO; digit3<=FIVE; end
      16'd5074: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ZERO; digit3<=FIVE; end
      16'd5075: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ZERO; digit3<=FIVE; end
      16'd5076: begin digit0<=SIX; digit1<=SEVEN; digit2<=ZERO; digit3<=FIVE; end
      16'd5077: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ZERO; digit3<=FIVE; end
      16'd5078: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ZERO; digit3<=FIVE; end
      16'd5079: begin digit0<=NINE; digit1<=SEVEN; digit2<=ZERO; digit3<=FIVE; end
      16'd5080: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ZERO; digit3<=FIVE; end
      16'd5081: begin digit0<=ONE; digit1<=EIGHT; digit2<=ZERO; digit3<=FIVE; end
      16'd5082: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ZERO; digit3<=FIVE; end
      16'd5083: begin digit0<=THREE; digit1<=EIGHT; digit2<=ZERO; digit3<=FIVE; end
      16'd5084: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ZERO; digit3<=FIVE; end
      16'd5085: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ZERO; digit3<=FIVE; end
      16'd5086: begin digit0<=SIX; digit1<=EIGHT; digit2<=ZERO; digit3<=FIVE; end
      16'd5087: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ZERO; digit3<=FIVE; end
      16'd5088: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ZERO; digit3<=FIVE; end
      16'd5089: begin digit0<=NINE; digit1<=EIGHT; digit2<=ZERO; digit3<=FIVE; end
      16'd5090: begin digit0<=ZERO; digit1<=NINE; digit2<=ZERO; digit3<=FIVE; end
      16'd5091: begin digit0<=ONE; digit1<=NINE; digit2<=ZERO; digit3<=FIVE; end
      16'd5092: begin digit0<=ZERO; digit1<=NINE; digit2<=ZERO; digit3<=FIVE; end
      16'd5093: begin digit0<=THREE; digit1<=NINE; digit2<=ZERO; digit3<=FIVE; end
      16'd5094: begin digit0<=FOUR; digit1<=NINE; digit2<=ZERO; digit3<=FIVE; end
      16'd5095: begin digit0<=FIVE; digit1<=NINE; digit2<=ZERO; digit3<=FIVE; end
      16'd5096: begin digit0<=SIX; digit1<=NINE; digit2<=ZERO; digit3<=FIVE; end
      16'd5097: begin digit0<=SEVEN; digit1<=NINE; digit2<=ZERO; digit3<=FIVE; end
      16'd5098: begin digit0<=EIGHT; digit1<=NINE; digit2<=ZERO; digit3<=FIVE; end
      16'd5099: begin digit0<=NINE; digit1<=NINE; digit2<=ZERO; digit3<=FIVE; end
	  16'd5100: begin digit0<=ZERO; digit1<=ZERO; digit2<=ONE; digit3<=FIVE; end
      16'd5101: begin digit0<=ONE; digit1<=ZERO; digit2<=ONE; digit3<=FIVE; end
      16'd5102: begin digit0<=TWO; digit1<=ZERO; digit2<=ONE; digit3<=FIVE; end
      16'd5103: begin digit0<=THREE; digit1<=ZERO; digit2<=ONE; digit3<=FIVE; end
      16'd5104: begin digit0<=FOUR; digit1<=ZERO; digit2<=ONE; digit3<=FIVE; end
      16'd5105: begin digit0<=FIVE; digit1<=ZERO; digit2<=ONE; digit3<=FIVE; end
      16'd5106: begin digit0<=SIX; digit1<=ZERO; digit2<=ONE; digit3<=FIVE; end
      16'd5107: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ONE; digit3<=FIVE; end
      16'd5108: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ONE; digit3<=FIVE; end
      16'd5109: begin digit0<=NINE; digit1<=ZERO; digit2<=ONE; digit3<=FIVE; end
      16'd5110: begin digit0<=ZERO; digit1<=ONE; digit2<=ONE; digit3<=FIVE; end
      16'd5111: begin digit0<=ONE; digit1<=ONE; digit2<=ONE; digit3<=FIVE; end
      16'd5112: begin digit0<=TWO; digit1<=ONE; digit2<=ONE; digit3<=FIVE; end
      16'd5113: begin digit0<=THREE; digit1<=ONE; digit2<=ONE; digit3<=FIVE; end
      16'd5114: begin digit0<=FOUR; digit1<=ONE; digit2<=ONE; digit3<=FIVE; end
      16'd5115: begin digit0<=FIVE; digit1<=ONE; digit2<=ONE; digit3<=FIVE; end
      16'd5116: begin digit0<=SIX; digit1<=ONE; digit2<=ONE; digit3<=FIVE; end
      16'd5117: begin digit0<=SEVEN; digit1<=ONE; digit2<=ONE; digit3<=FIVE; end
      16'd5118: begin digit0<=EIGHT; digit1<=ONE; digit2<=ONE; digit3<=FIVE; end
      16'd5119: begin digit0<=NINE; digit1<=ONE; digit2<=ONE; digit3<=FIVE; end
      16'd5120: begin digit0<=ZERO; digit1<=TWO; digit2<=ONE; digit3<=FIVE; end
      16'd5121: begin digit0<=ONE; digit1<=TWO; digit2<=ONE; digit3<=FIVE; end
      16'd5122: begin digit0<=TWO; digit1<=TWO; digit2<=ONE; digit3<=FIVE; end
      16'd5123: begin digit0<=THREE; digit1<=TWO; digit2<=ONE; digit3<=FIVE; end
      16'd5124: begin digit0<=FOUR; digit1<=TWO; digit2<=ONE; digit3<=FIVE; end
      16'd5125: begin digit0<=FIVE; digit1<=TWO; digit2<=ONE; digit3<=FIVE; end
      16'd5126: begin digit0<=SIX; digit1<=TWO; digit2<=ONE; digit3<=FIVE; end
      16'd5127: begin digit0<=SEVEN; digit1<=TWO; digit2<=ONE; digit3<=FIVE; end
      16'd5128: begin digit0<=EIGHT; digit1<=TWO; digit2<=ONE; digit3<=FIVE; end
      16'd5129: begin digit0<=NINE; digit1<=TWO; digit2<=ONE; digit3<=FIVE; end
      16'd5130: begin digit0<=ZERO; digit1<=THREE; digit2<=ONE; digit3<=FIVE; end
      16'd5131: begin digit0<=ONE; digit1<=THREE; digit2<=ONE; digit3<=FIVE; end
      16'd5132: begin digit0<=TWO; digit1<=THREE; digit2<=ONE; digit3<=FIVE; end
      16'd5133: begin digit0<=THREE; digit1<=THREE; digit2<=ONE; digit3<=FIVE; end
      16'd5134: begin digit0<=FOUR; digit1<=THREE; digit2<=ONE; digit3<=FIVE; end
      16'd5135: begin digit0<=FIVE; digit1<=THREE; digit2<=ONE; digit3<=FIVE; end
      16'd5136: begin digit0<=SIX; digit1<=THREE; digit2<=ONE; digit3<=FIVE; end
      16'd5137: begin digit0<=SEVEN; digit1<=THREE; digit2<=ONE; digit3<=FIVE; end
      16'd5138: begin digit0<=EIGHT; digit1<=THREE; digit2<=ONE; digit3<=FIVE; end
      16'd5139: begin digit0<=NINE; digit1<=THREE; digit2<=ONE; digit3<=FIVE; end
      16'd5140: begin digit0<=ZERO; digit1<=FOUR; digit2<=ONE; digit3<=FIVE; end
      16'd5141: begin digit0<=ONE; digit1<=FOUR; digit2<=ONE; digit3<=FIVE; end
      16'd5142: begin digit0<=TWO; digit1<=FOUR; digit2<=ONE; digit3<=FIVE; end
      16'd5143: begin digit0<=THREE; digit1<=FOUR; digit2<=ONE; digit3<=FIVE; end
      16'd5144: begin digit0<=FOUR; digit1<=FOUR; digit2<=ONE; digit3<=FIVE; end
      16'd5145: begin digit0<=FIVE; digit1<=FOUR; digit2<=ONE; digit3<=FIVE; end
      16'd5146: begin digit0<=SIX; digit1<=FOUR; digit2<=ONE; digit3<=FIVE; end
      16'd5147: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ONE; digit3<=FIVE; end
      16'd5148: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ONE; digit3<=FIVE; end
      16'd5149: begin digit0<=NINE; digit1<=FOUR; digit2<=ONE; digit3<=FIVE; end
      16'd5150: begin digit0<=ZERO; digit1<=FIVE; digit2<=ONE; digit3<=FIVE; end
      16'd5151: begin digit0<=ONE; digit1<=FIVE; digit2<=ONE; digit3<=FIVE; end
      16'd5152: begin digit0<=TWO; digit1<=FIVE; digit2<=ONE; digit3<=FIVE; end
      16'd5153: begin digit0<=THREE; digit1<=FIVE; digit2<=ONE; digit3<=FIVE; end
      16'd5154: begin digit0<=FOUR; digit1<=FIVE; digit2<=ONE; digit3<=FIVE; end
      16'd5155: begin digit0<=FIVE; digit1<=FIVE; digit2<=ONE; digit3<=FIVE; end
      16'd5156: begin digit0<=SIX; digit1<=FIVE; digit2<=ONE; digit3<=FIVE; end
      16'd5157: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ONE; digit3<=FIVE; end
      16'd5158: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ONE; digit3<=FIVE; end
      16'd5159: begin digit0<=NINE; digit1<=FIVE; digit2<=ONE; digit3<=FIVE; end
      16'd5160: begin digit0<=ZERO; digit1<=SIX; digit2<=ONE; digit3<=FIVE; end
      16'd5161: begin digit0<=ONE; digit1<=SIX; digit2<=ONE; digit3<=FIVE; end
      16'd5162: begin digit0<=TWO; digit1<=SIX; digit2<=ONE; digit3<=FIVE; end
      16'd5163: begin digit0<=THREE; digit1<=SIX; digit2<=ONE; digit3<=FIVE; end
      16'd5164: begin digit0<=FOUR; digit1<=SIX; digit2<=ONE; digit3<=FIVE; end
      16'd5165: begin digit0<=FIVE; digit1<=SIX; digit2<=ONE; digit3<=FIVE; end
      16'd5166: begin digit0<=SIX; digit1<=SIX; digit2<=ONE; digit3<=FIVE; end
      16'd5167: begin digit0<=SEVEN; digit1<=SIX; digit2<=ONE; digit3<=FIVE; end
      16'd5168: begin digit0<=EIGHT; digit1<=SIX; digit2<=ONE; digit3<=FIVE; end
      16'd5169: begin digit0<=NINE; digit1<=SIX; digit2<=ONE; digit3<=FIVE; end
      16'd5170: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ONE; digit3<=FIVE; end
      16'd5171: begin digit0<=ONE; digit1<=SEVEN; digit2<=ONE; digit3<=FIVE; end
      16'd5172: begin digit0<=TWO; digit1<=SEVEN; digit2<=ONE; digit3<=FIVE; end
      16'd5173: begin digit0<=THREE; digit1<=SEVEN; digit2<=ONE; digit3<=FIVE; end
      16'd5174: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ONE; digit3<=FIVE; end
      16'd5175: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ONE; digit3<=FIVE; end
      16'd5176: begin digit0<=SIX; digit1<=SEVEN; digit2<=ONE; digit3<=FIVE; end
      16'd5177: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ONE; digit3<=FIVE; end
      16'd5178: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ONE; digit3<=FIVE; end
      16'd5179: begin digit0<=NINE; digit1<=SEVEN; digit2<=ONE; digit3<=FIVE; end
      16'd5180: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=FIVE; end
      16'd5181: begin digit0<=ONE; digit1<=EIGHT; digit2<=ONE; digit3<=FIVE; end
      16'd5182: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=FIVE; end
      16'd5183: begin digit0<=THREE; digit1<=EIGHT; digit2<=ONE; digit3<=FIVE; end
      16'd5184: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ONE; digit3<=FIVE; end
      16'd5185: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ONE; digit3<=FIVE; end
      16'd5186: begin digit0<=SIX; digit1<=EIGHT; digit2<=ONE; digit3<=FIVE; end
      16'd5187: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ONE; digit3<=FIVE; end
      16'd5188: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ONE; digit3<=FIVE; end
      16'd5189: begin digit0<=NINE; digit1<=EIGHT; digit2<=ONE; digit3<=FIVE; end
      16'd5190: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=FIVE; end
      16'd5191: begin digit0<=ONE; digit1<=NINE; digit2<=ONE; digit3<=FIVE; end
      16'd5192: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=FIVE; end
      16'd5193: begin digit0<=THREE; digit1<=NINE; digit2<=ONE; digit3<=FIVE; end
      16'd5194: begin digit0<=FOUR; digit1<=NINE; digit2<=ONE; digit3<=FIVE; end
      16'd5195: begin digit0<=FIVE; digit1<=NINE; digit2<=ONE; digit3<=FIVE; end
      16'd5196: begin digit0<=SIX; digit1<=NINE; digit2<=ONE; digit3<=FIVE; end
      16'd5197: begin digit0<=SEVEN; digit1<=NINE; digit2<=ONE; digit3<=FIVE; end
      16'd5198: begin digit0<=EIGHT; digit1<=NINE; digit2<=ONE; digit3<=FIVE; end
      16'd5199: begin digit0<=NINE; digit1<=NINE; digit2<=ONE; digit3<=FIVE; end
	  16'd5200: begin digit0<=ZERO; digit1<=ZERO; digit2<=TWO; digit3<=FIVE; end
      16'd5201: begin digit0<=ONE; digit1<=ZERO; digit2<=TWO; digit3<=FIVE; end
      16'd5202: begin digit0<=TWO; digit1<=ZERO; digit2<=TWO; digit3<=FIVE; end
      16'd5203: begin digit0<=THREE; digit1<=ZERO; digit2<=TWO; digit3<=FIVE; end
      16'd5204: begin digit0<=FOUR; digit1<=ZERO; digit2<=TWO; digit3<=FIVE; end
      16'd5205: begin digit0<=FIVE; digit1<=ZERO; digit2<=TWO; digit3<=FIVE; end
      16'd5206: begin digit0<=SIX; digit1<=ZERO; digit2<=TWO; digit3<=FIVE; end
      16'd5207: begin digit0<=SEVEN; digit1<=ZERO; digit2<=TWO; digit3<=FIVE; end
      16'd5208: begin digit0<=EIGHT; digit1<=ZERO; digit2<=TWO; digit3<=FIVE; end
      16'd5209: begin digit0<=NINE; digit1<=ZERO; digit2<=TWO; digit3<=FIVE; end
      16'd5210: begin digit0<=ZERO; digit1<=ONE; digit2<=TWO; digit3<=FIVE; end
      16'd5211: begin digit0<=ONE; digit1<=ONE; digit2<=TWO; digit3<=FIVE; end
      16'd5212: begin digit0<=TWO; digit1<=ONE; digit2<=TWO; digit3<=FIVE; end
      16'd5213: begin digit0<=THREE; digit1<=ONE; digit2<=TWO; digit3<=FIVE; end
      16'd5214: begin digit0<=FOUR; digit1<=ONE; digit2<=TWO; digit3<=FIVE; end
      16'd5215: begin digit0<=FIVE; digit1<=ONE; digit2<=TWO; digit3<=FIVE; end
      16'd5216: begin digit0<=SIX; digit1<=ONE; digit2<=TWO; digit3<=FIVE; end
      16'd5217: begin digit0<=SEVEN; digit1<=ONE; digit2<=TWO; digit3<=FIVE; end
      16'd5218: begin digit0<=EIGHT; digit1<=ONE; digit2<=TWO; digit3<=FIVE; end
      16'd5219: begin digit0<=NINE; digit1<=ONE; digit2<=TWO; digit3<=FIVE; end
      16'd5220: begin digit0<=ZERO; digit1<=TWO; digit2<=TWO; digit3<=FIVE; end
      16'd5221: begin digit0<=ONE; digit1<=TWO; digit2<=TWO; digit3<=FIVE; end
      16'd5222: begin digit0<=TWO; digit1<=TWO; digit2<=TWO; digit3<=FIVE; end
      16'd5223: begin digit0<=THREE; digit1<=TWO; digit2<=TWO; digit3<=FIVE; end
      16'd5224: begin digit0<=FOUR; digit1<=TWO; digit2<=TWO; digit3<=FIVE; end
      16'd5225: begin digit0<=FIVE; digit1<=TWO; digit2<=TWO; digit3<=FIVE; end
      16'd5226: begin digit0<=SIX; digit1<=TWO; digit2<=TWO; digit3<=FIVE; end
      16'd5227: begin digit0<=SEVEN; digit1<=TWO; digit2<=TWO; digit3<=FIVE; end
      16'd5228: begin digit0<=EIGHT; digit1<=TWO; digit2<=TWO; digit3<=FIVE; end
      16'd5229: begin digit0<=NINE; digit1<=TWO; digit2<=TWO; digit3<=FIVE; end
      16'd5230: begin digit0<=ZERO; digit1<=THREE; digit2<=TWO; digit3<=FIVE; end
      16'd5231: begin digit0<=ONE; digit1<=THREE; digit2<=TWO; digit3<=FIVE; end
      16'd5232: begin digit0<=TWO; digit1<=THREE; digit2<=TWO; digit3<=FIVE; end
      16'd5233: begin digit0<=THREE; digit1<=THREE; digit2<=TWO; digit3<=FIVE; end
      16'd5234: begin digit0<=FOUR; digit1<=THREE; digit2<=TWO; digit3<=FIVE; end
      16'd5235: begin digit0<=FIVE; digit1<=THREE; digit2<=TWO; digit3<=FIVE; end
      16'd5236: begin digit0<=SIX; digit1<=THREE; digit2<=TWO; digit3<=FIVE; end
      16'd5237: begin digit0<=SEVEN; digit1<=THREE; digit2<=TWO; digit3<=FIVE; end
      16'd5238: begin digit0<=EIGHT; digit1<=THREE; digit2<=TWO; digit3<=FIVE; end
      16'd5239: begin digit0<=NINE; digit1<=THREE; digit2<=TWO; digit3<=FIVE; end
      16'd5240: begin digit0<=ZERO; digit1<=FOUR; digit2<=TWO; digit3<=FIVE; end
      16'd5241: begin digit0<=ONE; digit1<=FOUR; digit2<=TWO; digit3<=FIVE; end
      16'd5242: begin digit0<=TWO; digit1<=FOUR; digit2<=TWO; digit3<=FIVE; end
      16'd5243: begin digit0<=THREE; digit1<=FOUR; digit2<=TWO; digit3<=FIVE; end
      16'd5244: begin digit0<=FOUR; digit1<=FOUR; digit2<=TWO; digit3<=FIVE; end
      16'd5245: begin digit0<=FIVE; digit1<=FOUR; digit2<=TWO; digit3<=FIVE; end
      16'd5246: begin digit0<=SIX; digit1<=FOUR; digit2<=TWO; digit3<=FIVE; end
      16'd5247: begin digit0<=SEVEN; digit1<=FOUR; digit2<=TWO; digit3<=FIVE; end
      16'd5248: begin digit0<=EIGHT; digit1<=FOUR; digit2<=TWO; digit3<=FIVE; end
      16'd5249: begin digit0<=NINE; digit1<=FOUR; digit2<=TWO; digit3<=FIVE; end
      16'd5250: begin digit0<=ZERO; digit1<=FIVE; digit2<=TWO; digit3<=FIVE; end
      16'd5251: begin digit0<=ONE; digit1<=FIVE; digit2<=TWO; digit3<=FIVE; end
      16'd5252: begin digit0<=TWO; digit1<=FIVE; digit2<=TWO; digit3<=FIVE; end
      16'd5253: begin digit0<=THREE; digit1<=FIVE; digit2<=TWO; digit3<=FIVE; end
      16'd5254: begin digit0<=FOUR; digit1<=FIVE; digit2<=TWO; digit3<=FIVE; end
      16'd5255: begin digit0<=FIVE; digit1<=FIVE; digit2<=TWO; digit3<=FIVE; end
      16'd5256: begin digit0<=SIX; digit1<=FIVE; digit2<=TWO; digit3<=FIVE; end
      16'd5257: begin digit0<=SEVEN; digit1<=FIVE; digit2<=TWO; digit3<=FIVE; end
      16'd5258: begin digit0<=EIGHT; digit1<=FIVE; digit2<=TWO; digit3<=FIVE; end
      16'd5259: begin digit0<=NINE; digit1<=FIVE; digit2<=TWO; digit3<=FIVE; end
      16'd5260: begin digit0<=ZERO; digit1<=SIX; digit2<=TWO; digit3<=FIVE; end
      16'd5261: begin digit0<=ONE; digit1<=SIX; digit2<=TWO; digit3<=FIVE; end
      16'd5262: begin digit0<=TWO; digit1<=SIX; digit2<=TWO; digit3<=FIVE; end
      16'd5263: begin digit0<=THREE; digit1<=SIX; digit2<=TWO; digit3<=FIVE; end
      16'd5264: begin digit0<=FOUR; digit1<=SIX; digit2<=TWO; digit3<=FIVE; end
      16'd5265: begin digit0<=FIVE; digit1<=SIX; digit2<=TWO; digit3<=FIVE; end
      16'd5266: begin digit0<=SIX; digit1<=SIX; digit2<=TWO; digit3<=FIVE; end
      16'd5267: begin digit0<=SEVEN; digit1<=SIX; digit2<=TWO; digit3<=FIVE; end
      16'd5268: begin digit0<=EIGHT; digit1<=SIX; digit2<=TWO; digit3<=FIVE; end
      16'd5269: begin digit0<=NINE; digit1<=SIX; digit2<=TWO; digit3<=FIVE; end
      16'd5270: begin digit0<=ZERO; digit1<=SEVEN; digit2<=TWO; digit3<=FIVE; end
      16'd5271: begin digit0<=ONE; digit1<=SEVEN; digit2<=TWO; digit3<=FIVE; end
      16'd5272: begin digit0<=TWO; digit1<=SEVEN; digit2<=TWO; digit3<=FIVE; end
      16'd5273: begin digit0<=THREE; digit1<=SEVEN; digit2<=TWO; digit3<=FIVE; end
      16'd5274: begin digit0<=FOUR; digit1<=SEVEN; digit2<=TWO; digit3<=FIVE; end
      16'd5275: begin digit0<=FIVE; digit1<=SEVEN; digit2<=TWO; digit3<=FIVE; end
      16'd5276: begin digit0<=SIX; digit1<=SEVEN; digit2<=TWO; digit3<=FIVE; end
      16'd5277: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=TWO; digit3<=FIVE; end
      16'd5278: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=TWO; digit3<=FIVE; end
      16'd5279: begin digit0<=NINE; digit1<=SEVEN; digit2<=TWO; digit3<=FIVE; end
      16'd5280: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=FIVE; end
      16'd5281: begin digit0<=ONE; digit1<=EIGHT; digit2<=TWO; digit3<=FIVE; end
      16'd5282: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=FIVE; end
      16'd5283: begin digit0<=THREE; digit1<=EIGHT; digit2<=TWO; digit3<=FIVE; end
      16'd5284: begin digit0<=FOUR; digit1<=EIGHT; digit2<=TWO; digit3<=FIVE; end
      16'd5285: begin digit0<=FIVE; digit1<=EIGHT; digit2<=TWO; digit3<=FIVE; end
      16'd5286: begin digit0<=SIX; digit1<=EIGHT; digit2<=TWO; digit3<=FIVE; end
      16'd5287: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=TWO; digit3<=FIVE; end
      16'd5288: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=TWO; digit3<=FIVE; end
      16'd5289: begin digit0<=NINE; digit1<=EIGHT; digit2<=TWO; digit3<=FIVE; end
      16'd5290: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=FIVE; end
      16'd5291: begin digit0<=ONE; digit1<=NINE; digit2<=TWO; digit3<=FIVE; end
      16'd5292: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=FIVE; end
      16'd5293: begin digit0<=THREE; digit1<=NINE; digit2<=TWO; digit3<=FIVE; end
      16'd5294: begin digit0<=FOUR; digit1<=NINE; digit2<=TWO; digit3<=FIVE; end
      16'd5295: begin digit0<=FIVE; digit1<=NINE; digit2<=TWO; digit3<=FIVE; end
      16'd5296: begin digit0<=SIX; digit1<=NINE; digit2<=TWO; digit3<=FIVE; end
      16'd5297: begin digit0<=SEVEN; digit1<=NINE; digit2<=TWO; digit3<=FIVE; end
      16'd5298: begin digit0<=EIGHT; digit1<=NINE; digit2<=TWO; digit3<=FIVE; end
      16'd5299: begin digit0<=NINE; digit1<=NINE; digit2<=TWO; digit3<=FIVE; end
	  16'd5300: begin digit0<=ZERO; digit1<=ZERO; digit2<=THREE; digit3<=FIVE; end
      16'd5301: begin digit0<=ONE; digit1<=ZERO; digit2<=THREE; digit3<=FIVE; end
      16'd5302: begin digit0<=TWO; digit1<=ZERO; digit2<=THREE; digit3<=FIVE; end
      16'd5303: begin digit0<=THREE; digit1<=ZERO; digit2<=THREE; digit3<=FIVE; end
      16'd5304: begin digit0<=FOUR; digit1<=ZERO; digit2<=THREE; digit3<=FIVE; end
      16'd5305: begin digit0<=FIVE; digit1<=ZERO; digit2<=THREE; digit3<=FIVE; end
      16'd5306: begin digit0<=SIX; digit1<=ZERO; digit2<=THREE; digit3<=FIVE; end
      16'd5307: begin digit0<=SEVEN; digit1<=ZERO; digit2<=THREE; digit3<=FIVE; end
      16'd5308: begin digit0<=EIGHT; digit1<=ZERO; digit2<=THREE; digit3<=FIVE; end
      16'd5309: begin digit0<=NINE; digit1<=ZERO; digit2<=THREE; digit3<=FIVE; end
      16'd5310: begin digit0<=ZERO; digit1<=ONE; digit2<=THREE; digit3<=FIVE; end
      16'd5311: begin digit0<=ONE; digit1<=ONE; digit2<=THREE; digit3<=FIVE; end
      16'd5312: begin digit0<=TWO; digit1<=ONE; digit2<=THREE; digit3<=FIVE; end
      16'd5313: begin digit0<=THREE; digit1<=ONE; digit2<=THREE; digit3<=FIVE; end
      16'd5314: begin digit0<=FOUR; digit1<=ONE; digit2<=THREE; digit3<=FIVE; end
      16'd5315: begin digit0<=FIVE; digit1<=ONE; digit2<=THREE; digit3<=FIVE; end
      16'd5316: begin digit0<=SIX; digit1<=ONE; digit2<=THREE; digit3<=FIVE; end
      16'd5317: begin digit0<=SEVEN; digit1<=ONE; digit2<=THREE; digit3<=FIVE; end
      16'd5318: begin digit0<=EIGHT; digit1<=ONE; digit2<=THREE; digit3<=FIVE; end
      16'd5319: begin digit0<=NINE; digit1<=ONE; digit2<=THREE; digit3<=FIVE; end
      16'd5320: begin digit0<=ZERO; digit1<=TWO; digit2<=THREE; digit3<=FIVE; end
      16'd5321: begin digit0<=ONE; digit1<=TWO; digit2<=THREE; digit3<=FIVE; end
      16'd5322: begin digit0<=TWO; digit1<=TWO; digit2<=THREE; digit3<=FIVE; end
      16'd5323: begin digit0<=THREE; digit1<=TWO; digit2<=THREE; digit3<=FIVE; end
      16'd5324: begin digit0<=FOUR; digit1<=TWO; digit2<=THREE; digit3<=FIVE; end
      16'd5325: begin digit0<=FIVE; digit1<=TWO; digit2<=THREE; digit3<=FIVE; end
      16'd5326: begin digit0<=SIX; digit1<=TWO; digit2<=THREE; digit3<=FIVE; end
      16'd5327: begin digit0<=SEVEN; digit1<=TWO; digit2<=THREE; digit3<=FIVE; end
      16'd5328: begin digit0<=EIGHT; digit1<=TWO; digit2<=THREE; digit3<=FIVE; end
      16'd5329: begin digit0<=NINE; digit1<=TWO; digit2<=THREE; digit3<=FIVE; end
      16'd5330: begin digit0<=ZERO; digit1<=THREE; digit2<=THREE; digit3<=FIVE; end
      16'd5331: begin digit0<=ONE; digit1<=THREE; digit2<=THREE; digit3<=FIVE; end
      16'd5332: begin digit0<=TWO; digit1<=THREE; digit2<=THREE; digit3<=FIVE; end
      16'd5333: begin digit0<=THREE; digit1<=THREE; digit2<=THREE; digit3<=FIVE; end
      16'd5334: begin digit0<=FOUR; digit1<=THREE; digit2<=THREE; digit3<=FIVE; end
      16'd5335: begin digit0<=FIVE; digit1<=THREE; digit2<=THREE; digit3<=FIVE; end
      16'd5336: begin digit0<=SIX; digit1<=THREE; digit2<=THREE; digit3<=FIVE; end
      16'd5337: begin digit0<=SEVEN; digit1<=THREE; digit2<=THREE; digit3<=FIVE; end
      16'd5338: begin digit0<=EIGHT; digit1<=THREE; digit2<=THREE; digit3<=FIVE; end
      16'd5339: begin digit0<=NINE; digit1<=THREE; digit2<=THREE; digit3<=FIVE; end
      16'd5340: begin digit0<=ZERO; digit1<=FOUR; digit2<=THREE; digit3<=FIVE; end
      16'd5341: begin digit0<=ONE; digit1<=FOUR; digit2<=THREE; digit3<=FIVE; end
      16'd5342: begin digit0<=TWO; digit1<=FOUR; digit2<=THREE; digit3<=FIVE; end
      16'd5343: begin digit0<=THREE; digit1<=FOUR; digit2<=THREE; digit3<=FIVE; end
      16'd5344: begin digit0<=FOUR; digit1<=FOUR; digit2<=THREE; digit3<=FIVE; end
      16'd5345: begin digit0<=FIVE; digit1<=FOUR; digit2<=THREE; digit3<=FIVE; end
      16'd5346: begin digit0<=SIX; digit1<=FOUR; digit2<=THREE; digit3<=FIVE; end
      16'd5347: begin digit0<=SEVEN; digit1<=FOUR; digit2<=THREE; digit3<=FIVE; end
      16'd5348: begin digit0<=EIGHT; digit1<=FOUR; digit2<=THREE; digit3<=FIVE; end
      16'd5349: begin digit0<=NINE; digit1<=FOUR; digit2<=THREE; digit3<=FIVE; end
      16'd5350: begin digit0<=ZERO; digit1<=FIVE; digit2<=THREE; digit3<=FIVE; end
      16'd5351: begin digit0<=ONE; digit1<=FIVE; digit2<=THREE; digit3<=FIVE; end
      16'd5352: begin digit0<=TWO; digit1<=FIVE; digit2<=THREE; digit3<=FIVE; end
      16'd5353: begin digit0<=THREE; digit1<=FIVE; digit2<=THREE; digit3<=FIVE; end
      16'd5354: begin digit0<=FOUR; digit1<=FIVE; digit2<=THREE; digit3<=FIVE; end
      16'd5355: begin digit0<=FIVE; digit1<=FIVE; digit2<=THREE; digit3<=FIVE; end
      16'd5356: begin digit0<=SIX; digit1<=FIVE; digit2<=THREE; digit3<=FIVE; end
      16'd5357: begin digit0<=SEVEN; digit1<=FIVE; digit2<=THREE; digit3<=FIVE; end
      16'd5358: begin digit0<=EIGHT; digit1<=FIVE; digit2<=THREE; digit3<=FIVE; end
      16'd5359: begin digit0<=NINE; digit1<=FIVE; digit2<=THREE; digit3<=FIVE; end
      16'd5360: begin digit0<=ZERO; digit1<=SIX; digit2<=THREE; digit3<=FIVE; end
      16'd5361: begin digit0<=ONE; digit1<=SIX; digit2<=THREE; digit3<=FIVE; end
      16'd5362: begin digit0<=TWO; digit1<=SIX; digit2<=THREE; digit3<=FIVE; end
      16'd5363: begin digit0<=THREE; digit1<=SIX; digit2<=THREE; digit3<=FIVE; end
      16'd5364: begin digit0<=FOUR; digit1<=SIX; digit2<=THREE; digit3<=FIVE; end
      16'd5365: begin digit0<=FIVE; digit1<=SIX; digit2<=THREE; digit3<=FIVE; end
      16'd5366: begin digit0<=SIX; digit1<=SIX; digit2<=THREE; digit3<=FIVE; end
      16'd5367: begin digit0<=SEVEN; digit1<=SIX; digit2<=THREE; digit3<=FIVE; end
      16'd5368: begin digit0<=EIGHT; digit1<=SIX; digit2<=THREE; digit3<=FIVE; end
      16'd5369: begin digit0<=NINE; digit1<=SIX; digit2<=THREE; digit3<=FIVE; end
      16'd5370: begin digit0<=ZERO; digit1<=SEVEN; digit2<=THREE; digit3<=FIVE; end
      16'd5371: begin digit0<=ONE; digit1<=SEVEN; digit2<=THREE; digit3<=FIVE; end
      16'd5372: begin digit0<=TWO; digit1<=SEVEN; digit2<=THREE; digit3<=FIVE; end
      16'd5373: begin digit0<=THREE; digit1<=SEVEN; digit2<=THREE; digit3<=FIVE; end
      16'd5374: begin digit0<=FOUR; digit1<=SEVEN; digit2<=THREE; digit3<=FIVE; end
      16'd5375: begin digit0<=FIVE; digit1<=SEVEN; digit2<=THREE; digit3<=FIVE; end
      16'd5376: begin digit0<=SIX; digit1<=SEVEN; digit2<=THREE; digit3<=FIVE; end
      16'd5377: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=THREE; digit3<=FIVE; end
      16'd5378: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=THREE; digit3<=FIVE; end
      16'd5379: begin digit0<=NINE; digit1<=SEVEN; digit2<=THREE; digit3<=FIVE; end
      16'd5380: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=FIVE; end
      16'd5381: begin digit0<=ONE; digit1<=EIGHT; digit2<=THREE; digit3<=FIVE; end
      16'd5382: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=FIVE; end
      16'd5383: begin digit0<=THREE; digit1<=EIGHT; digit2<=THREE; digit3<=FIVE; end
      16'd5384: begin digit0<=FOUR; digit1<=EIGHT; digit2<=THREE; digit3<=FIVE; end
      16'd5385: begin digit0<=FIVE; digit1<=EIGHT; digit2<=THREE; digit3<=FIVE; end
      16'd5386: begin digit0<=SIX; digit1<=EIGHT; digit2<=THREE; digit3<=FIVE; end
      16'd5387: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=THREE; digit3<=FIVE; end
      16'd5388: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=THREE; digit3<=FIVE; end
      16'd5389: begin digit0<=NINE; digit1<=EIGHT; digit2<=THREE; digit3<=FIVE; end
      16'd5390: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=FIVE; end
      16'd5391: begin digit0<=ONE; digit1<=NINE; digit2<=THREE; digit3<=FIVE; end
      16'd5392: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=FIVE; end
      16'd5393: begin digit0<=THREE; digit1<=NINE; digit2<=THREE; digit3<=FIVE; end
      16'd5394: begin digit0<=FOUR; digit1<=NINE; digit2<=THREE; digit3<=FIVE; end
      16'd5395: begin digit0<=FIVE; digit1<=NINE; digit2<=THREE; digit3<=FIVE; end
      16'd5396: begin digit0<=SIX; digit1<=NINE; digit2<=THREE; digit3<=FIVE; end
      16'd5397: begin digit0<=SEVEN; digit1<=NINE; digit2<=THREE; digit3<=FIVE; end
      16'd5398: begin digit0<=EIGHT; digit1<=NINE; digit2<=THREE; digit3<=FIVE; end
      16'd5399: begin digit0<=NINE; digit1<=NINE; digit2<=THREE; digit3<=FIVE; end
	  16'd5400: begin digit0<=ZERO; digit1<=ZERO; digit2<=FOUR; digit3<=FIVE; end
      16'd5401: begin digit0<=ONE; digit1<=ZERO; digit2<=FOUR; digit3<=FIVE; end
      16'd5402: begin digit0<=TWO; digit1<=ZERO; digit2<=FOUR; digit3<=FIVE; end
      16'd5403: begin digit0<=THREE; digit1<=ZERO; digit2<=FOUR; digit3<=FIVE; end
      16'd5404: begin digit0<=FOUR; digit1<=ZERO; digit2<=FOUR; digit3<=FIVE; end
      16'd5405: begin digit0<=FIVE; digit1<=ZERO; digit2<=FOUR; digit3<=FIVE; end
      16'd5406: begin digit0<=SIX; digit1<=ZERO; digit2<=FOUR; digit3<=FIVE; end
      16'd5407: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FOUR; digit3<=FIVE; end
      16'd5408: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FOUR; digit3<=FIVE; end
      16'd5409: begin digit0<=NINE; digit1<=ZERO; digit2<=FOUR; digit3<=FIVE; end
      16'd5410: begin digit0<=ZERO; digit1<=ONE; digit2<=FOUR; digit3<=FIVE; end
      16'd5411: begin digit0<=ONE; digit1<=ONE; digit2<=FOUR; digit3<=FIVE; end
      16'd5412: begin digit0<=TWO; digit1<=ONE; digit2<=FOUR; digit3<=FIVE; end
      16'd5413: begin digit0<=THREE; digit1<=ONE; digit2<=FOUR; digit3<=FIVE; end
      16'd5414: begin digit0<=FOUR; digit1<=ONE; digit2<=FOUR; digit3<=FIVE; end
      16'd5415: begin digit0<=FIVE; digit1<=ONE; digit2<=FOUR; digit3<=FIVE; end
      16'd5416: begin digit0<=SIX; digit1<=ONE; digit2<=FOUR; digit3<=FIVE; end
      16'd5417: begin digit0<=SEVEN; digit1<=ONE; digit2<=FOUR; digit3<=FIVE; end
      16'd5418: begin digit0<=EIGHT; digit1<=ONE; digit2<=FOUR; digit3<=FIVE; end
      16'd5419: begin digit0<=NINE; digit1<=ONE; digit2<=FOUR; digit3<=FIVE; end
      16'd5420: begin digit0<=ZERO; digit1<=TWO; digit2<=FOUR; digit3<=FIVE; end
      16'd5421: begin digit0<=ONE; digit1<=TWO; digit2<=FOUR; digit3<=FIVE; end
      16'd5422: begin digit0<=TWO; digit1<=TWO; digit2<=FOUR; digit3<=FIVE; end
      16'd5423: begin digit0<=THREE; digit1<=TWO; digit2<=FOUR; digit3<=FIVE; end
      16'd5424: begin digit0<=FOUR; digit1<=TWO; digit2<=FOUR; digit3<=FIVE; end
      16'd5425: begin digit0<=FIVE; digit1<=TWO; digit2<=FOUR; digit3<=FIVE; end
      16'd5426: begin digit0<=SIX; digit1<=TWO; digit2<=FOUR; digit3<=FIVE; end
      16'd5427: begin digit0<=SEVEN; digit1<=TWO; digit2<=FOUR; digit3<=FIVE; end
      16'd5428: begin digit0<=EIGHT; digit1<=TWO; digit2<=FOUR; digit3<=FIVE; end
      16'd5429: begin digit0<=NINE; digit1<=TWO; digit2<=FOUR; digit3<=FIVE; end
      16'd5430: begin digit0<=ZERO; digit1<=THREE; digit2<=FOUR; digit3<=FIVE; end
      16'd5431: begin digit0<=ONE; digit1<=THREE; digit2<=FOUR; digit3<=FIVE; end
      16'd5432: begin digit0<=TWO; digit1<=THREE; digit2<=FOUR; digit3<=FIVE; end
      16'd5433: begin digit0<=THREE; digit1<=THREE; digit2<=FOUR; digit3<=FIVE; end
      16'd5434: begin digit0<=FOUR; digit1<=THREE; digit2<=FOUR; digit3<=FIVE; end
      16'd5435: begin digit0<=FIVE; digit1<=THREE; digit2<=FOUR; digit3<=FIVE; end
      16'd5436: begin digit0<=SIX; digit1<=THREE; digit2<=FOUR; digit3<=FIVE; end
      16'd5437: begin digit0<=SEVEN; digit1<=THREE; digit2<=FOUR; digit3<=FIVE; end
      16'd5438: begin digit0<=EIGHT; digit1<=THREE; digit2<=FOUR; digit3<=FIVE; end
      16'd5439: begin digit0<=NINE; digit1<=THREE; digit2<=FOUR; digit3<=FIVE; end
      16'd5440: begin digit0<=ZERO; digit1<=FOUR; digit2<=FOUR; digit3<=FIVE; end
      16'd5441: begin digit0<=ONE; digit1<=FOUR; digit2<=FOUR; digit3<=FIVE; end
      16'd5442: begin digit0<=TWO; digit1<=FOUR; digit2<=FOUR; digit3<=FIVE; end
      16'd5443: begin digit0<=THREE; digit1<=FOUR; digit2<=FOUR; digit3<=FIVE; end
      16'd5444: begin digit0<=FOUR; digit1<=FOUR; digit2<=FOUR; digit3<=FIVE; end
      16'd5445: begin digit0<=FIVE; digit1<=FOUR; digit2<=FOUR; digit3<=FIVE; end
      16'd5446: begin digit0<=SIX; digit1<=FOUR; digit2<=FOUR; digit3<=FIVE; end
      16'd5447: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FOUR; digit3<=FIVE; end
      16'd5448: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FOUR; digit3<=FIVE; end
      16'd5449: begin digit0<=NINE; digit1<=FOUR; digit2<=FOUR; digit3<=FIVE; end
      16'd5450: begin digit0<=ZERO; digit1<=FIVE; digit2<=FOUR; digit3<=FIVE; end
      16'd5451: begin digit0<=ONE; digit1<=FIVE; digit2<=FOUR; digit3<=FIVE; end
      16'd5452: begin digit0<=TWO; digit1<=FIVE; digit2<=FOUR; digit3<=FIVE; end
      16'd5453: begin digit0<=THREE; digit1<=FIVE; digit2<=FOUR; digit3<=FIVE; end
      16'd5454: begin digit0<=FOUR; digit1<=FIVE; digit2<=FOUR; digit3<=FIVE; end
      16'd5455: begin digit0<=FIVE; digit1<=FIVE; digit2<=FOUR; digit3<=FIVE; end
      16'd5456: begin digit0<=SIX; digit1<=FIVE; digit2<=FOUR; digit3<=FIVE; end
      16'd5457: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FOUR; digit3<=FIVE; end
      16'd5458: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FOUR; digit3<=FIVE; end
      16'd5459: begin digit0<=NINE; digit1<=FIVE; digit2<=FOUR; digit3<=FIVE; end
      16'd5460: begin digit0<=ZERO; digit1<=SIX; digit2<=FOUR; digit3<=FIVE; end
      16'd5461: begin digit0<=ONE; digit1<=SIX; digit2<=FOUR; digit3<=FIVE; end
      16'd5462: begin digit0<=TWO; digit1<=SIX; digit2<=FOUR; digit3<=FIVE; end
      16'd5463: begin digit0<=THREE; digit1<=SIX; digit2<=FOUR; digit3<=FIVE; end
      16'd5464: begin digit0<=FOUR; digit1<=SIX; digit2<=FOUR; digit3<=FIVE; end
      16'd5465: begin digit0<=FIVE; digit1<=SIX; digit2<=FOUR; digit3<=FIVE; end
      16'd5466: begin digit0<=SIX; digit1<=SIX; digit2<=FOUR; digit3<=FIVE; end
      16'd5467: begin digit0<=SEVEN; digit1<=SIX; digit2<=FOUR; digit3<=FIVE; end
      16'd5468: begin digit0<=EIGHT; digit1<=SIX; digit2<=FOUR; digit3<=FIVE; end
      16'd5469: begin digit0<=NINE; digit1<=SIX; digit2<=FOUR; digit3<=FIVE; end
      16'd5470: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FOUR; digit3<=FIVE; end
      16'd5471: begin digit0<=ONE; digit1<=SEVEN; digit2<=FOUR; digit3<=FIVE; end
      16'd5472: begin digit0<=TWO; digit1<=SEVEN; digit2<=FOUR; digit3<=FIVE; end
      16'd5473: begin digit0<=THREE; digit1<=SEVEN; digit2<=FOUR; digit3<=FIVE; end
      16'd5474: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FOUR; digit3<=FIVE; end
      16'd5475: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FOUR; digit3<=FIVE; end
      16'd5476: begin digit0<=SIX; digit1<=SEVEN; digit2<=FOUR; digit3<=FIVE; end
      16'd5477: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FOUR; digit3<=FIVE; end
      16'd5478: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FOUR; digit3<=FIVE; end
      16'd5479: begin digit0<=NINE; digit1<=SEVEN; digit2<=FOUR; digit3<=FIVE; end
      16'd5480: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=FIVE; end
      16'd5481: begin digit0<=ONE; digit1<=EIGHT; digit2<=FOUR; digit3<=FIVE; end
      16'd5482: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=FIVE; end
      16'd5483: begin digit0<=THREE; digit1<=EIGHT; digit2<=FOUR; digit3<=FIVE; end
      16'd5484: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FOUR; digit3<=FIVE; end
      16'd5485: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FOUR; digit3<=FIVE; end
      16'd5486: begin digit0<=SIX; digit1<=EIGHT; digit2<=FOUR; digit3<=FIVE; end
      16'd5487: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FOUR; digit3<=FIVE; end
      16'd5488: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FOUR; digit3<=FIVE; end
      16'd5489: begin digit0<=NINE; digit1<=EIGHT; digit2<=FOUR; digit3<=FIVE; end
      16'd5490: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=FIVE; end
      16'd5491: begin digit0<=ONE; digit1<=NINE; digit2<=FOUR; digit3<=FIVE; end
      16'd5492: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=FIVE; end
      16'd5493: begin digit0<=THREE; digit1<=NINE; digit2<=FOUR; digit3<=FIVE; end
      16'd5494: begin digit0<=FOUR; digit1<=NINE; digit2<=FOUR; digit3<=FIVE; end
      16'd5495: begin digit0<=FIVE; digit1<=NINE; digit2<=FOUR; digit3<=FIVE; end
      16'd5496: begin digit0<=SIX; digit1<=NINE; digit2<=FOUR; digit3<=FIVE; end
      16'd5497: begin digit0<=SEVEN; digit1<=NINE; digit2<=FOUR; digit3<=FIVE; end
      16'd5498: begin digit0<=EIGHT; digit1<=NINE; digit2<=FOUR; digit3<=FIVE; end
      16'd5499: begin digit0<=NINE; digit1<=NINE; digit2<=FOUR; digit3<=FIVE; end
	  16'd5500: begin digit0<=ZERO; digit1<=ZERO; digit2<=FIVE; digit3<=FIVE; end
      16'd5501: begin digit0<=ONE; digit1<=ZERO; digit2<=FIVE; digit3<=FIVE; end
      16'd5502: begin digit0<=TWO; digit1<=ZERO; digit2<=FIVE; digit3<=FIVE; end
      16'd5503: begin digit0<=THREE; digit1<=ZERO; digit2<=FIVE; digit3<=FIVE; end
      16'd5504: begin digit0<=FOUR; digit1<=ZERO; digit2<=FIVE; digit3<=FIVE; end
      16'd5505: begin digit0<=FIVE; digit1<=ZERO; digit2<=FIVE; digit3<=FIVE; end
      16'd5506: begin digit0<=SIX; digit1<=ZERO; digit2<=FIVE; digit3<=FIVE; end
      16'd5507: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FIVE; digit3<=FIVE; end
      16'd5508: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FIVE; digit3<=FIVE; end
      16'd5509: begin digit0<=NINE; digit1<=ZERO; digit2<=FIVE; digit3<=FIVE; end
      16'd5510: begin digit0<=ZERO; digit1<=ONE; digit2<=FIVE; digit3<=FIVE; end
      16'd5511: begin digit0<=ONE; digit1<=ONE; digit2<=FIVE; digit3<=FIVE; end
      16'd5512: begin digit0<=TWO; digit1<=ONE; digit2<=FIVE; digit3<=FIVE; end
      16'd5513: begin digit0<=THREE; digit1<=ONE; digit2<=FIVE; digit3<=FIVE; end
      16'd5514: begin digit0<=FOUR; digit1<=ONE; digit2<=FIVE; digit3<=FIVE; end
      16'd5515: begin digit0<=FIVE; digit1<=ONE; digit2<=FIVE; digit3<=FIVE; end
      16'd5516: begin digit0<=SIX; digit1<=ONE; digit2<=FIVE; digit3<=FIVE; end
      16'd5517: begin digit0<=SEVEN; digit1<=ONE; digit2<=FIVE; digit3<=FIVE; end
      16'd5518: begin digit0<=EIGHT; digit1<=ONE; digit2<=FIVE; digit3<=FIVE; end
      16'd5519: begin digit0<=NINE; digit1<=ONE; digit2<=FIVE; digit3<=FIVE; end
      16'd5520: begin digit0<=ZERO; digit1<=TWO; digit2<=FIVE; digit3<=FIVE; end
      16'd5521: begin digit0<=ONE; digit1<=TWO; digit2<=FIVE; digit3<=FIVE; end
      16'd5522: begin digit0<=TWO; digit1<=TWO; digit2<=FIVE; digit3<=FIVE; end
      16'd5523: begin digit0<=THREE; digit1<=TWO; digit2<=FIVE; digit3<=FIVE; end
      16'd5524: begin digit0<=FOUR; digit1<=TWO; digit2<=FIVE; digit3<=FIVE; end
      16'd5525: begin digit0<=FIVE; digit1<=TWO; digit2<=FIVE; digit3<=FIVE; end
      16'd5526: begin digit0<=SIX; digit1<=TWO; digit2<=FIVE; digit3<=FIVE; end
      16'd5527: begin digit0<=SEVEN; digit1<=TWO; digit2<=FIVE; digit3<=FIVE; end
      16'd5528: begin digit0<=EIGHT; digit1<=TWO; digit2<=FIVE; digit3<=FIVE; end
      16'd5529: begin digit0<=NINE; digit1<=TWO; digit2<=FIVE; digit3<=FIVE; end
      16'd5530: begin digit0<=ZERO; digit1<=THREE; digit2<=FIVE; digit3<=FIVE; end
      16'd5531: begin digit0<=ONE; digit1<=THREE; digit2<=FIVE; digit3<=FIVE; end
      16'd5532: begin digit0<=TWO; digit1<=THREE; digit2<=FIVE; digit3<=FIVE; end
      16'd5533: begin digit0<=THREE; digit1<=THREE; digit2<=FIVE; digit3<=FIVE; end
      16'd5534: begin digit0<=FOUR; digit1<=THREE; digit2<=FIVE; digit3<=FIVE; end
      16'd5535: begin digit0<=FIVE; digit1<=THREE; digit2<=FIVE; digit3<=FIVE; end
      16'd5536: begin digit0<=SIX; digit1<=THREE; digit2<=FIVE; digit3<=FIVE; end
      16'd5537: begin digit0<=SEVEN; digit1<=THREE; digit2<=FIVE; digit3<=FIVE; end
      16'd5538: begin digit0<=EIGHT; digit1<=THREE; digit2<=FIVE; digit3<=FIVE; end
      16'd5539: begin digit0<=NINE; digit1<=THREE; digit2<=FIVE; digit3<=FIVE; end
      16'd5540: begin digit0<=ZERO; digit1<=FOUR; digit2<=FIVE; digit3<=FIVE; end
      16'd5541: begin digit0<=ONE; digit1<=FOUR; digit2<=FIVE; digit3<=FIVE; end
      16'd5542: begin digit0<=TWO; digit1<=FOUR; digit2<=FIVE; digit3<=FIVE; end
      16'd5543: begin digit0<=THREE; digit1<=FOUR; digit2<=FIVE; digit3<=FIVE; end
      16'd5544: begin digit0<=FOUR; digit1<=FOUR; digit2<=FIVE; digit3<=FIVE; end
      16'd5545: begin digit0<=FIVE; digit1<=FOUR; digit2<=FIVE; digit3<=FIVE; end
      16'd5546: begin digit0<=SIX; digit1<=FOUR; digit2<=FIVE; digit3<=FIVE; end
      16'd5547: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FIVE; digit3<=FIVE; end
      16'd5548: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FIVE; digit3<=FIVE; end
      16'd5549: begin digit0<=NINE; digit1<=FOUR; digit2<=FIVE; digit3<=FIVE; end
      16'd5550: begin digit0<=ZERO; digit1<=FIVE; digit2<=FIVE; digit3<=FIVE; end
      16'd5551: begin digit0<=ONE; digit1<=FIVE; digit2<=FIVE; digit3<=FIVE; end
      16'd5552: begin digit0<=TWO; digit1<=FIVE; digit2<=FIVE; digit3<=FIVE; end
      16'd5553: begin digit0<=THREE; digit1<=FIVE; digit2<=FIVE; digit3<=FIVE; end
      16'd5554: begin digit0<=FOUR; digit1<=FIVE; digit2<=FIVE; digit3<=FIVE; end
      16'd5555: begin digit0<=FIVE; digit1<=FIVE; digit2<=FIVE; digit3<=FIVE; end
      16'd5556: begin digit0<=SIX; digit1<=FIVE; digit2<=FIVE; digit3<=FIVE; end
      16'd5557: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FIVE; digit3<=FIVE; end
      16'd5558: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FIVE; digit3<=FIVE; end
      16'd5559: begin digit0<=NINE; digit1<=FIVE; digit2<=FIVE; digit3<=FIVE; end
      16'd5560: begin digit0<=ZERO; digit1<=SIX; digit2<=FIVE; digit3<=FIVE; end
      16'd5561: begin digit0<=ONE; digit1<=SIX; digit2<=FIVE; digit3<=FIVE; end
      16'd5562: begin digit0<=TWO; digit1<=SIX; digit2<=FIVE; digit3<=FIVE; end
      16'd5563: begin digit0<=THREE; digit1<=SIX; digit2<=FIVE; digit3<=FIVE; end
      16'd5564: begin digit0<=FOUR; digit1<=SIX; digit2<=FIVE; digit3<=FIVE; end
      16'd5565: begin digit0<=FIVE; digit1<=SIX; digit2<=FIVE; digit3<=FIVE; end
      16'd5566: begin digit0<=SIX; digit1<=SIX; digit2<=FIVE; digit3<=FIVE; end
      16'd5567: begin digit0<=SEVEN; digit1<=SIX; digit2<=FIVE; digit3<=FIVE; end
      16'd5568: begin digit0<=EIGHT; digit1<=SIX; digit2<=FIVE; digit3<=FIVE; end
      16'd5569: begin digit0<=NINE; digit1<=SIX; digit2<=FIVE; digit3<=FIVE; end
      16'd5570: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FIVE; digit3<=FIVE; end
      16'd5571: begin digit0<=ONE; digit1<=SEVEN; digit2<=FIVE; digit3<=FIVE; end
      16'd5572: begin digit0<=TWO; digit1<=SEVEN; digit2<=FIVE; digit3<=FIVE; end
      16'd5573: begin digit0<=THREE; digit1<=SEVEN; digit2<=FIVE; digit3<=FIVE; end
      16'd5574: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FIVE; digit3<=FIVE; end
      16'd5575: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FIVE; digit3<=FIVE; end
      16'd5576: begin digit0<=SIX; digit1<=SEVEN; digit2<=FIVE; digit3<=FIVE; end
      16'd5577: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FIVE; digit3<=FIVE; end
      16'd5578: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FIVE; digit3<=FIVE; end
      16'd5579: begin digit0<=NINE; digit1<=SEVEN; digit2<=FIVE; digit3<=FIVE; end
      16'd5580: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=FIVE; end
      16'd5581: begin digit0<=ONE; digit1<=EIGHT; digit2<=FIVE; digit3<=FIVE; end
      16'd5582: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=FIVE; end
      16'd5583: begin digit0<=THREE; digit1<=EIGHT; digit2<=FIVE; digit3<=FIVE; end
      16'd5584: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FIVE; digit3<=FIVE; end
      16'd5585: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FIVE; digit3<=FIVE; end
      16'd5586: begin digit0<=SIX; digit1<=EIGHT; digit2<=FIVE; digit3<=FIVE; end
      16'd5587: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FIVE; digit3<=FIVE; end
      16'd5588: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FIVE; digit3<=FIVE; end
      16'd5589: begin digit0<=NINE; digit1<=EIGHT; digit2<=FIVE; digit3<=FIVE; end
      16'd5590: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=FIVE; end
      16'd5591: begin digit0<=ONE; digit1<=NINE; digit2<=FIVE; digit3<=FIVE; end
      16'd5592: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=FIVE; end
      16'd5593: begin digit0<=THREE; digit1<=NINE; digit2<=FIVE; digit3<=FIVE; end
      16'd5594: begin digit0<=FOUR; digit1<=NINE; digit2<=FIVE; digit3<=FIVE; end
      16'd5595: begin digit0<=FIVE; digit1<=NINE; digit2<=FIVE; digit3<=FIVE; end
      16'd5596: begin digit0<=SIX; digit1<=NINE; digit2<=FIVE; digit3<=FIVE; end
      16'd5597: begin digit0<=SEVEN; digit1<=NINE; digit2<=FIVE; digit3<=FIVE; end
      16'd5598: begin digit0<=EIGHT; digit1<=NINE; digit2<=FIVE; digit3<=FIVE; end
      16'd5599: begin digit0<=NINE; digit1<=NINE; digit2<=FIVE; digit3<=FIVE; end
	  16'd5600: begin digit0<=ZERO; digit1<=ZERO; digit2<=SIX; digit3<=FIVE; end
      16'd5601: begin digit0<=ONE; digit1<=ZERO; digit2<=SIX; digit3<=FIVE; end
      16'd5602: begin digit0<=TWO; digit1<=ZERO; digit2<=SIX; digit3<=FIVE; end
      16'd5603: begin digit0<=THREE; digit1<=ZERO; digit2<=SIX; digit3<=FIVE; end
      16'd5604: begin digit0<=FOUR; digit1<=ZERO; digit2<=SIX; digit3<=FIVE; end
      16'd5605: begin digit0<=FIVE; digit1<=ZERO; digit2<=SIX; digit3<=FIVE; end
      16'd5606: begin digit0<=SIX; digit1<=ZERO; digit2<=SIX; digit3<=FIVE; end
      16'd5607: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SIX; digit3<=FIVE; end
      16'd5608: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SIX; digit3<=FIVE; end
      16'd5609: begin digit0<=NINE; digit1<=ZERO; digit2<=SIX; digit3<=FIVE; end
      16'd5610: begin digit0<=ZERO; digit1<=ONE; digit2<=SIX; digit3<=FIVE; end
      16'd5611: begin digit0<=ONE; digit1<=ONE; digit2<=SIX; digit3<=FIVE; end
      16'd5612: begin digit0<=TWO; digit1<=ONE; digit2<=SIX; digit3<=FIVE; end
      16'd5613: begin digit0<=THREE; digit1<=ONE; digit2<=SIX; digit3<=FIVE; end
      16'd5614: begin digit0<=FOUR; digit1<=ONE; digit2<=SIX; digit3<=FIVE; end
      16'd5615: begin digit0<=FIVE; digit1<=ONE; digit2<=SIX; digit3<=FIVE; end
      16'd5616: begin digit0<=SIX; digit1<=ONE; digit2<=SIX; digit3<=FIVE; end
      16'd5617: begin digit0<=SEVEN; digit1<=ONE; digit2<=SIX; digit3<=FIVE; end
      16'd5618: begin digit0<=EIGHT; digit1<=ONE; digit2<=SIX; digit3<=FIVE; end
      16'd5619: begin digit0<=NINE; digit1<=ONE; digit2<=SIX; digit3<=FIVE; end
      16'd5620: begin digit0<=ZERO; digit1<=TWO; digit2<=SIX; digit3<=FIVE; end
      16'd5621: begin digit0<=ONE; digit1<=TWO; digit2<=SIX; digit3<=FIVE; end
      16'd5622: begin digit0<=TWO; digit1<=TWO; digit2<=SIX; digit3<=FIVE; end
      16'd5623: begin digit0<=THREE; digit1<=TWO; digit2<=SIX; digit3<=FIVE; end
      16'd5624: begin digit0<=FOUR; digit1<=TWO; digit2<=SIX; digit3<=FIVE; end
      16'd5625: begin digit0<=FIVE; digit1<=TWO; digit2<=SIX; digit3<=FIVE; end
      16'd5626: begin digit0<=SIX; digit1<=TWO; digit2<=SIX; digit3<=FIVE; end
      16'd5627: begin digit0<=SEVEN; digit1<=TWO; digit2<=SIX; digit3<=FIVE; end
      16'd5628: begin digit0<=EIGHT; digit1<=TWO; digit2<=SIX; digit3<=FIVE; end
      16'd5629: begin digit0<=NINE; digit1<=TWO; digit2<=SIX; digit3<=FIVE; end
      16'd5630: begin digit0<=ZERO; digit1<=THREE; digit2<=SIX; digit3<=FIVE; end
      16'd5631: begin digit0<=ONE; digit1<=THREE; digit2<=SIX; digit3<=FIVE; end
      16'd5632: begin digit0<=TWO; digit1<=THREE; digit2<=SIX; digit3<=FIVE; end
      16'd5633: begin digit0<=THREE; digit1<=THREE; digit2<=SIX; digit3<=FIVE; end
      16'd5634: begin digit0<=FOUR; digit1<=THREE; digit2<=SIX; digit3<=FIVE; end
      16'd5635: begin digit0<=FIVE; digit1<=THREE; digit2<=SIX; digit3<=FIVE; end
      16'd5636: begin digit0<=SIX; digit1<=THREE; digit2<=SIX; digit3<=FIVE; end
      16'd5637: begin digit0<=SEVEN; digit1<=THREE; digit2<=SIX; digit3<=FIVE; end
      16'd5638: begin digit0<=EIGHT; digit1<=THREE; digit2<=SIX; digit3<=FIVE; end
      16'd5639: begin digit0<=NINE; digit1<=THREE; digit2<=SIX; digit3<=FIVE; end
      16'd5640: begin digit0<=ZERO; digit1<=FOUR; digit2<=SIX; digit3<=FIVE; end
      16'd5641: begin digit0<=ONE; digit1<=FOUR; digit2<=SIX; digit3<=FIVE; end
      16'd5642: begin digit0<=TWO; digit1<=FOUR; digit2<=SIX; digit3<=FIVE; end
      16'd5643: begin digit0<=THREE; digit1<=FOUR; digit2<=SIX; digit3<=FIVE; end
      16'd5644: begin digit0<=FOUR; digit1<=FOUR; digit2<=SIX; digit3<=FIVE; end
      16'd5645: begin digit0<=FIVE; digit1<=FOUR; digit2<=SIX; digit3<=FIVE; end
      16'd5646: begin digit0<=SIX; digit1<=FOUR; digit2<=SIX; digit3<=FIVE; end
      16'd5647: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SIX; digit3<=FIVE; end
      16'd5648: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SIX; digit3<=FIVE; end
      16'd5649: begin digit0<=NINE; digit1<=FOUR; digit2<=SIX; digit3<=FIVE; end
      16'd5650: begin digit0<=ZERO; digit1<=FIVE; digit2<=SIX; digit3<=FIVE; end
      16'd5651: begin digit0<=ONE; digit1<=FIVE; digit2<=SIX; digit3<=FIVE; end
      16'd5652: begin digit0<=TWO; digit1<=FIVE; digit2<=SIX; digit3<=FIVE; end
      16'd5653: begin digit0<=THREE; digit1<=FIVE; digit2<=SIX; digit3<=FIVE; end
      16'd5654: begin digit0<=FOUR; digit1<=FIVE; digit2<=SIX; digit3<=FIVE; end
      16'd5655: begin digit0<=FIVE; digit1<=FIVE; digit2<=SIX; digit3<=FIVE; end
      16'd5656: begin digit0<=SIX; digit1<=FIVE; digit2<=SIX; digit3<=FIVE; end
      16'd5657: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SIX; digit3<=FIVE; end
      16'd5658: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SIX; digit3<=FIVE; end
      16'd5659: begin digit0<=NINE; digit1<=FIVE; digit2<=SIX; digit3<=FIVE; end
      16'd5660: begin digit0<=ZERO; digit1<=SIX; digit2<=SIX; digit3<=FIVE; end
      16'd5661: begin digit0<=ONE; digit1<=SIX; digit2<=SIX; digit3<=FIVE; end
      16'd5662: begin digit0<=TWO; digit1<=SIX; digit2<=SIX; digit3<=FIVE; end
      16'd5663: begin digit0<=THREE; digit1<=SIX; digit2<=SIX; digit3<=FIVE; end
      16'd5664: begin digit0<=FOUR; digit1<=SIX; digit2<=SIX; digit3<=FIVE; end
      16'd5665: begin digit0<=FIVE; digit1<=SIX; digit2<=SIX; digit3<=FIVE; end
      16'd5666: begin digit0<=SIX; digit1<=SIX; digit2<=SIX; digit3<=FIVE; end
      16'd5667: begin digit0<=SEVEN; digit1<=SIX; digit2<=SIX; digit3<=FIVE; end
      16'd5668: begin digit0<=EIGHT; digit1<=SIX; digit2<=SIX; digit3<=FIVE; end
      16'd5669: begin digit0<=NINE; digit1<=SIX; digit2<=SIX; digit3<=FIVE; end
      16'd5670: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SIX; digit3<=FIVE; end
      16'd5671: begin digit0<=ONE; digit1<=SEVEN; digit2<=SIX; digit3<=FIVE; end
      16'd5672: begin digit0<=TWO; digit1<=SEVEN; digit2<=SIX; digit3<=FIVE; end
      16'd5673: begin digit0<=THREE; digit1<=SEVEN; digit2<=SIX; digit3<=FIVE; end
      16'd5674: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SIX; digit3<=FIVE; end
      16'd5675: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SIX; digit3<=FIVE; end
      16'd5676: begin digit0<=SIX; digit1<=SEVEN; digit2<=SIX; digit3<=FIVE; end
      16'd5677: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SIX; digit3<=FIVE; end
      16'd5678: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SIX; digit3<=FIVE; end
      16'd5679: begin digit0<=NINE; digit1<=SEVEN; digit2<=SIX; digit3<=FIVE; end
      16'd5680: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=FIVE; end
      16'd5681: begin digit0<=ONE; digit1<=EIGHT; digit2<=SIX; digit3<=FIVE; end
      16'd5682: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=FIVE; end
      16'd5683: begin digit0<=THREE; digit1<=EIGHT; digit2<=SIX; digit3<=FIVE; end
      16'd5684: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SIX; digit3<=FIVE; end
      16'd5685: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SIX; digit3<=FIVE; end
      16'd5686: begin digit0<=SIX; digit1<=EIGHT; digit2<=SIX; digit3<=FIVE; end
      16'd5687: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SIX; digit3<=FIVE; end
      16'd5688: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SIX; digit3<=FIVE; end
      16'd5689: begin digit0<=NINE; digit1<=EIGHT; digit2<=SIX; digit3<=FIVE; end
      16'd5690: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=FIVE; end
      16'd5691: begin digit0<=ONE; digit1<=NINE; digit2<=SIX; digit3<=FIVE; end
      16'd5692: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=FIVE; end
      16'd5693: begin digit0<=THREE; digit1<=NINE; digit2<=SIX; digit3<=FIVE; end
      16'd5694: begin digit0<=FOUR; digit1<=NINE; digit2<=SIX; digit3<=FIVE; end
      16'd5695: begin digit0<=FIVE; digit1<=NINE; digit2<=SIX; digit3<=FIVE; end
      16'd5696: begin digit0<=SIX; digit1<=NINE; digit2<=SIX; digit3<=FIVE; end
      16'd5697: begin digit0<=SEVEN; digit1<=NINE; digit2<=SIX; digit3<=FIVE; end
      16'd5698: begin digit0<=EIGHT; digit1<=NINE; digit2<=SIX; digit3<=FIVE; end
      16'd5699: begin digit0<=NINE; digit1<=NINE; digit2<=SIX; digit3<=FIVE; end
	  16'd5700: begin digit0<=ZERO; digit1<=ZERO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5701: begin digit0<=ONE; digit1<=ZERO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5702: begin digit0<=TWO; digit1<=ZERO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5703: begin digit0<=THREE; digit1<=ZERO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5704: begin digit0<=FOUR; digit1<=ZERO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5705: begin digit0<=FIVE; digit1<=ZERO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5706: begin digit0<=SIX; digit1<=ZERO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5707: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5708: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5709: begin digit0<=NINE; digit1<=ZERO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5710: begin digit0<=ZERO; digit1<=ONE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5711: begin digit0<=ONE; digit1<=ONE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5712: begin digit0<=TWO; digit1<=ONE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5713: begin digit0<=THREE; digit1<=ONE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5714: begin digit0<=FOUR; digit1<=ONE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5715: begin digit0<=FIVE; digit1<=ONE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5716: begin digit0<=SIX; digit1<=ONE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5717: begin digit0<=SEVEN; digit1<=ONE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5718: begin digit0<=EIGHT; digit1<=ONE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5719: begin digit0<=NINE; digit1<=ONE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5720: begin digit0<=ZERO; digit1<=TWO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5721: begin digit0<=ONE; digit1<=TWO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5722: begin digit0<=TWO; digit1<=TWO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5723: begin digit0<=THREE; digit1<=TWO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5724: begin digit0<=FOUR; digit1<=TWO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5725: begin digit0<=FIVE; digit1<=TWO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5726: begin digit0<=SIX; digit1<=TWO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5727: begin digit0<=SEVEN; digit1<=TWO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5728: begin digit0<=EIGHT; digit1<=TWO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5729: begin digit0<=NINE; digit1<=TWO; digit2<=SEVEN; digit3<=FIVE; end
      16'd5730: begin digit0<=ZERO; digit1<=THREE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5731: begin digit0<=ONE; digit1<=THREE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5732: begin digit0<=TWO; digit1<=THREE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5733: begin digit0<=THREE; digit1<=THREE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5734: begin digit0<=FOUR; digit1<=THREE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5735: begin digit0<=FIVE; digit1<=THREE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5736: begin digit0<=SIX; digit1<=THREE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5737: begin digit0<=SEVEN; digit1<=THREE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5738: begin digit0<=EIGHT; digit1<=THREE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5739: begin digit0<=NINE; digit1<=THREE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5740: begin digit0<=ZERO; digit1<=FOUR; digit2<=SEVEN; digit3<=FIVE; end
      16'd5741: begin digit0<=ONE; digit1<=FOUR; digit2<=SEVEN; digit3<=FIVE; end
      16'd5742: begin digit0<=TWO; digit1<=FOUR; digit2<=SEVEN; digit3<=FIVE; end
      16'd5743: begin digit0<=THREE; digit1<=FOUR; digit2<=SEVEN; digit3<=FIVE; end
      16'd5744: begin digit0<=FOUR; digit1<=FOUR; digit2<=SEVEN; digit3<=FIVE; end
      16'd5745: begin digit0<=FIVE; digit1<=FOUR; digit2<=SEVEN; digit3<=FIVE; end
      16'd5746: begin digit0<=SIX; digit1<=FOUR; digit2<=SEVEN; digit3<=FIVE; end
      16'd5747: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SEVEN; digit3<=FIVE; end
      16'd5748: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SEVEN; digit3<=FIVE; end
      16'd5749: begin digit0<=NINE; digit1<=FOUR; digit2<=SEVEN; digit3<=FIVE; end
      16'd5750: begin digit0<=ZERO; digit1<=FIVE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5751: begin digit0<=ONE; digit1<=FIVE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5752: begin digit0<=TWO; digit1<=FIVE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5753: begin digit0<=THREE; digit1<=FIVE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5754: begin digit0<=FOUR; digit1<=FIVE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5755: begin digit0<=FIVE; digit1<=FIVE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5756: begin digit0<=SIX; digit1<=FIVE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5757: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5758: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5759: begin digit0<=NINE; digit1<=FIVE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5760: begin digit0<=ZERO; digit1<=SIX; digit2<=SEVEN; digit3<=FIVE; end
      16'd5761: begin digit0<=ONE; digit1<=SIX; digit2<=SEVEN; digit3<=FIVE; end
      16'd5762: begin digit0<=TWO; digit1<=SIX; digit2<=SEVEN; digit3<=FIVE; end
      16'd5763: begin digit0<=THREE; digit1<=SIX; digit2<=SEVEN; digit3<=FIVE; end
      16'd5764: begin digit0<=FOUR; digit1<=SIX; digit2<=SEVEN; digit3<=FIVE; end
      16'd5765: begin digit0<=FIVE; digit1<=SIX; digit2<=SEVEN; digit3<=FIVE; end
      16'd5766: begin digit0<=SIX; digit1<=SIX; digit2<=SEVEN; digit3<=FIVE; end
      16'd5767: begin digit0<=SEVEN; digit1<=SIX; digit2<=SEVEN; digit3<=FIVE; end
      16'd5768: begin digit0<=EIGHT; digit1<=SIX; digit2<=SEVEN; digit3<=FIVE; end
      16'd5769: begin digit0<=NINE; digit1<=SIX; digit2<=SEVEN; digit3<=FIVE; end
      16'd5770: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SEVEN; digit3<=FIVE; end
      16'd5771: begin digit0<=ONE; digit1<=SEVEN; digit2<=SEVEN; digit3<=FIVE; end
      16'd5772: begin digit0<=TWO; digit1<=SEVEN; digit2<=SEVEN; digit3<=FIVE; end
      16'd5773: begin digit0<=THREE; digit1<=SEVEN; digit2<=SEVEN; digit3<=FIVE; end
      16'd5774: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SEVEN; digit3<=FIVE; end
      16'd5775: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SEVEN; digit3<=FIVE; end
      16'd5776: begin digit0<=SIX; digit1<=SEVEN; digit2<=SEVEN; digit3<=FIVE; end
      16'd5777: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SEVEN; digit3<=FIVE; end
      16'd5778: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SEVEN; digit3<=FIVE; end
      16'd5779: begin digit0<=NINE; digit1<=SEVEN; digit2<=SEVEN; digit3<=FIVE; end
      16'd5780: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=FIVE; end
      16'd5781: begin digit0<=ONE; digit1<=EIGHT; digit2<=SEVEN; digit3<=FIVE; end
      16'd5782: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=FIVE; end
      16'd5783: begin digit0<=THREE; digit1<=EIGHT; digit2<=SEVEN; digit3<=FIVE; end
      16'd5784: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SEVEN; digit3<=FIVE; end
      16'd5785: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SEVEN; digit3<=FIVE; end
      16'd5786: begin digit0<=SIX; digit1<=EIGHT; digit2<=SEVEN; digit3<=FIVE; end
      16'd5787: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SEVEN; digit3<=FIVE; end
      16'd5788: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SEVEN; digit3<=FIVE; end
      16'd5789: begin digit0<=NINE; digit1<=EIGHT; digit2<=SEVEN; digit3<=FIVE; end
      16'd5790: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5791: begin digit0<=ONE; digit1<=NINE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5792: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5793: begin digit0<=THREE; digit1<=NINE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5794: begin digit0<=FOUR; digit1<=NINE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5795: begin digit0<=FIVE; digit1<=NINE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5796: begin digit0<=SIX; digit1<=NINE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5797: begin digit0<=SEVEN; digit1<=NINE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5798: begin digit0<=EIGHT; digit1<=NINE; digit2<=SEVEN; digit3<=FIVE; end
      16'd5799: begin digit0<=NINE; digit1<=NINE; digit2<=SEVEN; digit3<=FIVE; end
	  16'd5800: begin digit0<=ZERO; digit1<=ZERO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5801: begin digit0<=ONE; digit1<=ZERO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5802: begin digit0<=TWO; digit1<=ZERO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5803: begin digit0<=THREE; digit1<=ZERO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5804: begin digit0<=FOUR; digit1<=ZERO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5805: begin digit0<=FIVE; digit1<=ZERO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5806: begin digit0<=SIX; digit1<=ZERO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5807: begin digit0<=SEVEN; digit1<=ZERO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5808: begin digit0<=EIGHT; digit1<=ZERO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5809: begin digit0<=NINE; digit1<=ZERO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5810: begin digit0<=ZERO; digit1<=ONE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5811: begin digit0<=ONE; digit1<=ONE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5812: begin digit0<=TWO; digit1<=ONE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5813: begin digit0<=THREE; digit1<=ONE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5814: begin digit0<=FOUR; digit1<=ONE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5815: begin digit0<=FIVE; digit1<=ONE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5816: begin digit0<=SIX; digit1<=ONE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5817: begin digit0<=SEVEN; digit1<=ONE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5818: begin digit0<=EIGHT; digit1<=ONE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5819: begin digit0<=NINE; digit1<=ONE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5820: begin digit0<=ZERO; digit1<=TWO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5821: begin digit0<=ONE; digit1<=TWO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5822: begin digit0<=TWO; digit1<=TWO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5823: begin digit0<=THREE; digit1<=TWO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5824: begin digit0<=FOUR; digit1<=TWO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5825: begin digit0<=FIVE; digit1<=TWO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5826: begin digit0<=SIX; digit1<=TWO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5827: begin digit0<=SEVEN; digit1<=TWO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5828: begin digit0<=EIGHT; digit1<=TWO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5829: begin digit0<=NINE; digit1<=TWO; digit2<=EIGHT; digit3<=FIVE; end
      16'd5830: begin digit0<=ZERO; digit1<=THREE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5831: begin digit0<=ONE; digit1<=THREE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5832: begin digit0<=TWO; digit1<=THREE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5833: begin digit0<=THREE; digit1<=THREE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5834: begin digit0<=FOUR; digit1<=THREE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5835: begin digit0<=FIVE; digit1<=THREE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5836: begin digit0<=SIX; digit1<=THREE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5837: begin digit0<=SEVEN; digit1<=THREE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5838: begin digit0<=EIGHT; digit1<=THREE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5839: begin digit0<=NINE; digit1<=THREE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5840: begin digit0<=ZERO; digit1<=FOUR; digit2<=EIGHT; digit3<=FIVE; end
      16'd5841: begin digit0<=ONE; digit1<=FOUR; digit2<=EIGHT; digit3<=FIVE; end
      16'd5842: begin digit0<=TWO; digit1<=FOUR; digit2<=EIGHT; digit3<=FIVE; end
      16'd5843: begin digit0<=THREE; digit1<=FOUR; digit2<=EIGHT; digit3<=FIVE; end
      16'd5844: begin digit0<=FOUR; digit1<=FOUR; digit2<=EIGHT; digit3<=FIVE; end
      16'd5845: begin digit0<=FIVE; digit1<=FOUR; digit2<=EIGHT; digit3<=FIVE; end
      16'd5846: begin digit0<=SIX; digit1<=FOUR; digit2<=EIGHT; digit3<=FIVE; end
      16'd5847: begin digit0<=SEVEN; digit1<=FOUR; digit2<=EIGHT; digit3<=FIVE; end
      16'd5848: begin digit0<=EIGHT; digit1<=FOUR; digit2<=EIGHT; digit3<=FIVE; end
      16'd5849: begin digit0<=NINE; digit1<=FOUR; digit2<=EIGHT; digit3<=FIVE; end
      16'd5850: begin digit0<=ZERO; digit1<=FIVE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5851: begin digit0<=ONE; digit1<=FIVE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5852: begin digit0<=TWO; digit1<=FIVE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5853: begin digit0<=THREE; digit1<=FIVE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5854: begin digit0<=FOUR; digit1<=FIVE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5855: begin digit0<=FIVE; digit1<=FIVE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5856: begin digit0<=SIX; digit1<=FIVE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5857: begin digit0<=SEVEN; digit1<=FIVE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5858: begin digit0<=EIGHT; digit1<=FIVE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5859: begin digit0<=NINE; digit1<=FIVE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5860: begin digit0<=ZERO; digit1<=SIX; digit2<=EIGHT; digit3<=FIVE; end
      16'd5861: begin digit0<=ONE; digit1<=SIX; digit2<=EIGHT; digit3<=FIVE; end
      16'd5862: begin digit0<=TWO; digit1<=SIX; digit2<=EIGHT; digit3<=FIVE; end
      16'd5863: begin digit0<=THREE; digit1<=SIX; digit2<=EIGHT; digit3<=FIVE; end
      16'd5864: begin digit0<=FOUR; digit1<=SIX; digit2<=EIGHT; digit3<=FIVE; end
      16'd5865: begin digit0<=FIVE; digit1<=SIX; digit2<=EIGHT; digit3<=FIVE; end
      16'd5866: begin digit0<=SIX; digit1<=SIX; digit2<=EIGHT; digit3<=FIVE; end
      16'd5867: begin digit0<=SEVEN; digit1<=SIX; digit2<=EIGHT; digit3<=FIVE; end
      16'd5868: begin digit0<=EIGHT; digit1<=SIX; digit2<=EIGHT; digit3<=FIVE; end
      16'd5869: begin digit0<=NINE; digit1<=SIX; digit2<=EIGHT; digit3<=FIVE; end
      16'd5870: begin digit0<=ZERO; digit1<=SEVEN; digit2<=EIGHT; digit3<=FIVE; end
      16'd5871: begin digit0<=ONE; digit1<=SEVEN; digit2<=EIGHT; digit3<=FIVE; end
      16'd5872: begin digit0<=TWO; digit1<=SEVEN; digit2<=EIGHT; digit3<=FIVE; end
      16'd5873: begin digit0<=THREE; digit1<=SEVEN; digit2<=EIGHT; digit3<=FIVE; end
      16'd5874: begin digit0<=FOUR; digit1<=SEVEN; digit2<=EIGHT; digit3<=FIVE; end
      16'd5875: begin digit0<=FIVE; digit1<=SEVEN; digit2<=EIGHT; digit3<=FIVE; end
      16'd5876: begin digit0<=SIX; digit1<=SEVEN; digit2<=EIGHT; digit3<=FIVE; end
      16'd5877: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=EIGHT; digit3<=FIVE; end
      16'd5878: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=EIGHT; digit3<=FIVE; end
      16'd5879: begin digit0<=NINE; digit1<=SEVEN; digit2<=EIGHT; digit3<=FIVE; end
      16'd5880: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=FIVE; end
      16'd5881: begin digit0<=ONE; digit1<=EIGHT; digit2<=EIGHT; digit3<=FIVE; end
      16'd5882: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=FIVE; end
      16'd5883: begin digit0<=THREE; digit1<=EIGHT; digit2<=EIGHT; digit3<=FIVE; end
      16'd5884: begin digit0<=FOUR; digit1<=EIGHT; digit2<=EIGHT; digit3<=FIVE; end
      16'd5885: begin digit0<=FIVE; digit1<=EIGHT; digit2<=EIGHT; digit3<=FIVE; end
      16'd5886: begin digit0<=SIX; digit1<=EIGHT; digit2<=EIGHT; digit3<=FIVE; end
      16'd5887: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=EIGHT; digit3<=FIVE; end
      16'd5888: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=EIGHT; digit3<=FIVE; end
      16'd5889: begin digit0<=NINE; digit1<=EIGHT; digit2<=EIGHT; digit3<=FIVE; end
      16'd5890: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5891: begin digit0<=ONE; digit1<=NINE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5892: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5893: begin digit0<=THREE; digit1<=NINE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5894: begin digit0<=FOUR; digit1<=NINE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5895: begin digit0<=FIVE; digit1<=NINE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5896: begin digit0<=SIX; digit1<=NINE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5897: begin digit0<=SEVEN; digit1<=NINE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5898: begin digit0<=EIGHT; digit1<=NINE; digit2<=EIGHT; digit3<=FIVE; end
      16'd5899: begin digit0<=NINE; digit1<=NINE; digit2<=EIGHT; digit3<=FIVE; end
	  16'd5900: begin digit0<=ZERO; digit1<=ZERO; digit2<=NINE; digit3<=FIVE; end
      16'd5901: begin digit0<=ONE; digit1<=ZERO; digit2<=NINE; digit3<=FIVE; end
      16'd5902: begin digit0<=TWO; digit1<=ZERO; digit2<=NINE; digit3<=FIVE; end
      16'd5903: begin digit0<=THREE; digit1<=ZERO; digit2<=NINE; digit3<=FIVE; end
      16'd5904: begin digit0<=FOUR; digit1<=ZERO; digit2<=NINE; digit3<=FIVE; end
      16'd5905: begin digit0<=FIVE; digit1<=ZERO; digit2<=NINE; digit3<=FIVE; end
      16'd5906: begin digit0<=SIX; digit1<=ZERO; digit2<=NINE; digit3<=FIVE; end
      16'd5907: begin digit0<=SEVEN; digit1<=ZERO; digit2<=NINE; digit3<=FIVE; end
      16'd5908: begin digit0<=EIGHT; digit1<=ZERO; digit2<=NINE; digit3<=FIVE; end
      16'd5909: begin digit0<=NINE; digit1<=ZERO; digit2<=NINE; digit3<=FIVE; end
      16'd5910: begin digit0<=ZERO; digit1<=ONE; digit2<=NINE; digit3<=FIVE; end
      16'd5911: begin digit0<=ONE; digit1<=ONE; digit2<=NINE; digit3<=FIVE; end
      16'd5912: begin digit0<=TWO; digit1<=ONE; digit2<=NINE; digit3<=FIVE; end
      16'd5913: begin digit0<=THREE; digit1<=ONE; digit2<=NINE; digit3<=FIVE; end
      16'd5914: begin digit0<=FOUR; digit1<=ONE; digit2<=NINE; digit3<=FIVE; end
      16'd5915: begin digit0<=FIVE; digit1<=ONE; digit2<=NINE; digit3<=FIVE; end
      16'd5916: begin digit0<=SIX; digit1<=ONE; digit2<=NINE; digit3<=FIVE; end
      16'd5917: begin digit0<=SEVEN; digit1<=ONE; digit2<=NINE; digit3<=FIVE; end
      16'd5918: begin digit0<=EIGHT; digit1<=ONE; digit2<=NINE; digit3<=FIVE; end
      16'd5919: begin digit0<=NINE; digit1<=ONE; digit2<=NINE; digit3<=FIVE; end
      16'd5920: begin digit0<=ZERO; digit1<=TWO; digit2<=NINE; digit3<=FIVE; end
      16'd5921: begin digit0<=ONE; digit1<=TWO; digit2<=NINE; digit3<=FIVE; end
      16'd5922: begin digit0<=TWO; digit1<=TWO; digit2<=NINE; digit3<=FIVE; end
      16'd5923: begin digit0<=THREE; digit1<=TWO; digit2<=NINE; digit3<=FIVE; end
      16'd5924: begin digit0<=FOUR; digit1<=TWO; digit2<=NINE; digit3<=FIVE; end
      16'd5925: begin digit0<=FIVE; digit1<=TWO; digit2<=NINE; digit3<=FIVE; end
      16'd5926: begin digit0<=SIX; digit1<=TWO; digit2<=NINE; digit3<=FIVE; end
      16'd5927: begin digit0<=SEVEN; digit1<=TWO; digit2<=NINE; digit3<=FIVE; end
      16'd5928: begin digit0<=EIGHT; digit1<=TWO; digit2<=NINE; digit3<=FIVE; end
      16'd5929: begin digit0<=NINE; digit1<=TWO; digit2<=NINE; digit3<=FIVE; end
      16'd5930: begin digit0<=ZERO; digit1<=THREE; digit2<=NINE; digit3<=FIVE; end
      16'd5931: begin digit0<=ONE; digit1<=THREE; digit2<=NINE; digit3<=FIVE; end
      16'd5932: begin digit0<=TWO; digit1<=THREE; digit2<=NINE; digit3<=FIVE; end
      16'd5933: begin digit0<=THREE; digit1<=THREE; digit2<=NINE; digit3<=FIVE; end
      16'd5934: begin digit0<=FOUR; digit1<=THREE; digit2<=NINE; digit3<=FIVE; end
      16'd5935: begin digit0<=FIVE; digit1<=THREE; digit2<=NINE; digit3<=FIVE; end
      16'd5936: begin digit0<=SIX; digit1<=THREE; digit2<=NINE; digit3<=FIVE; end
      16'd5937: begin digit0<=SEVEN; digit1<=THREE; digit2<=NINE; digit3<=FIVE; end
      16'd5938: begin digit0<=EIGHT; digit1<=THREE; digit2<=NINE; digit3<=FIVE; end
      16'd5939: begin digit0<=NINE; digit1<=THREE; digit2<=NINE; digit3<=FIVE; end
      16'd5940: begin digit0<=ZERO; digit1<=FOUR; digit2<=NINE; digit3<=FIVE; end
      16'd5941: begin digit0<=ONE; digit1<=FOUR; digit2<=NINE; digit3<=FIVE; end
      16'd5942: begin digit0<=TWO; digit1<=FOUR; digit2<=NINE; digit3<=FIVE; end
      16'd5943: begin digit0<=THREE; digit1<=FOUR; digit2<=NINE; digit3<=FIVE; end
      16'd5944: begin digit0<=FOUR; digit1<=FOUR; digit2<=NINE; digit3<=FIVE; end
      16'd5945: begin digit0<=FIVE; digit1<=FOUR; digit2<=NINE; digit3<=FIVE; end
      16'd5946: begin digit0<=SIX; digit1<=FOUR; digit2<=NINE; digit3<=FIVE; end
      16'd5947: begin digit0<=SEVEN; digit1<=FOUR; digit2<=NINE; digit3<=FIVE; end
      16'd5948: begin digit0<=EIGHT; digit1<=FOUR; digit2<=NINE; digit3<=FIVE; end
      16'd5949: begin digit0<=NINE; digit1<=FOUR; digit2<=NINE; digit3<=FIVE; end
      16'd5950: begin digit0<=ZERO; digit1<=FIVE; digit2<=NINE; digit3<=FIVE; end
      16'd5951: begin digit0<=ONE; digit1<=FIVE; digit2<=NINE; digit3<=FIVE; end
      16'd5952: begin digit0<=TWO; digit1<=FIVE; digit2<=NINE; digit3<=FIVE; end
      16'd5953: begin digit0<=THREE; digit1<=FIVE; digit2<=NINE; digit3<=FIVE; end
      16'd5954: begin digit0<=FOUR; digit1<=FIVE; digit2<=NINE; digit3<=FIVE; end
      16'd5955: begin digit0<=FIVE; digit1<=FIVE; digit2<=NINE; digit3<=FIVE; end
      16'd5956: begin digit0<=SIX; digit1<=FIVE; digit2<=NINE; digit3<=FIVE; end
      16'd5957: begin digit0<=SEVEN; digit1<=FIVE; digit2<=NINE; digit3<=FIVE; end
      16'd5958: begin digit0<=EIGHT; digit1<=FIVE; digit2<=NINE; digit3<=FIVE; end
      16'd5959: begin digit0<=NINE; digit1<=FIVE; digit2<=NINE; digit3<=FIVE; end
      16'd5960: begin digit0<=ZERO; digit1<=SIX; digit2<=NINE; digit3<=FIVE; end
      16'd5961: begin digit0<=ONE; digit1<=SIX; digit2<=NINE; digit3<=FIVE; end
      16'd5962: begin digit0<=TWO; digit1<=SIX; digit2<=NINE; digit3<=FIVE; end
      16'd5963: begin digit0<=THREE; digit1<=SIX; digit2<=NINE; digit3<=FIVE; end
      16'd5964: begin digit0<=FOUR; digit1<=SIX; digit2<=NINE; digit3<=FIVE; end
      16'd5965: begin digit0<=FIVE; digit1<=SIX; digit2<=NINE; digit3<=FIVE; end
      16'd5966: begin digit0<=SIX; digit1<=SIX; digit2<=NINE; digit3<=FIVE; end
      16'd5967: begin digit0<=SEVEN; digit1<=SIX; digit2<=NINE; digit3<=FIVE; end
      16'd5968: begin digit0<=EIGHT; digit1<=SIX; digit2<=NINE; digit3<=FIVE; end
      16'd5969: begin digit0<=NINE; digit1<=SIX; digit2<=NINE; digit3<=FIVE; end
      16'd5970: begin digit0<=ZERO; digit1<=SEVEN; digit2<=NINE; digit3<=FIVE; end
      16'd5971: begin digit0<=ONE; digit1<=SEVEN; digit2<=NINE; digit3<=FIVE; end
      16'd5972: begin digit0<=TWO; digit1<=SEVEN; digit2<=NINE; digit3<=FIVE; end
      16'd5973: begin digit0<=THREE; digit1<=SEVEN; digit2<=NINE; digit3<=FIVE; end
      16'd5974: begin digit0<=FOUR; digit1<=SEVEN; digit2<=NINE; digit3<=FIVE; end
      16'd5975: begin digit0<=FIVE; digit1<=SEVEN; digit2<=NINE; digit3<=FIVE; end
      16'd5976: begin digit0<=SIX; digit1<=SEVEN; digit2<=NINE; digit3<=FIVE; end
      16'd5977: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=NINE; digit3<=FIVE; end
      16'd5978: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=NINE; digit3<=FIVE; end
      16'd5979: begin digit0<=NINE; digit1<=SEVEN; digit2<=NINE; digit3<=FIVE; end
      16'd5980: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=FIVE; end
      16'd5981: begin digit0<=ONE; digit1<=EIGHT; digit2<=NINE; digit3<=FIVE; end
      16'd5982: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=FIVE; end
      16'd5983: begin digit0<=THREE; digit1<=EIGHT; digit2<=NINE; digit3<=FIVE; end
      16'd5984: begin digit0<=FOUR; digit1<=EIGHT; digit2<=NINE; digit3<=FIVE; end
      16'd5985: begin digit0<=FIVE; digit1<=EIGHT; digit2<=NINE; digit3<=FIVE; end
      16'd5986: begin digit0<=SIX; digit1<=EIGHT; digit2<=NINE; digit3<=FIVE; end
      16'd5987: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=NINE; digit3<=FIVE; end
      16'd5988: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=NINE; digit3<=FIVE; end
      16'd5989: begin digit0<=NINE; digit1<=EIGHT; digit2<=NINE; digit3<=FIVE; end
      16'd5990: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=FIVE; end
      16'd5991: begin digit0<=ONE; digit1<=NINE; digit2<=NINE; digit3<=FIVE; end
      16'd5992: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=FIVE; end
      16'd5993: begin digit0<=THREE; digit1<=NINE; digit2<=NINE; digit3<=FIVE; end
      16'd5994: begin digit0<=FOUR; digit1<=NINE; digit2<=NINE; digit3<=FIVE; end
      16'd5995: begin digit0<=FIVE; digit1<=NINE; digit2<=NINE; digit3<=FIVE; end
      16'd5996: begin digit0<=SIX; digit1<=NINE; digit2<=NINE; digit3<=FIVE; end
      16'd5997: begin digit0<=SEVEN; digit1<=NINE; digit2<=NINE; digit3<=FIVE; end
      16'd5998: begin digit0<=EIGHT; digit1<=NINE; digit2<=NINE; digit3<=FIVE; end
      16'd5999: begin digit0<=NINE; digit1<=NINE; digit2<=NINE; digit3<=FIVE; end
	  16'd6000: begin digit0<=ZERO; digit1<=ZERO; digit2<=ZERO; digit3<=SIX; end
      16'd6001: begin digit0<=ONE; digit1<=ZERO; digit2<=ZERO; digit3<=SIX; end
      16'd6002: begin digit0<=TWO; digit1<=ZERO; digit2<=ZERO; digit3<=SIX; end
      16'd6003: begin digit0<=THREE; digit1<=ZERO; digit2<=ZERO; digit3<=SIX; end
      16'd6004: begin digit0<=FOUR; digit1<=ZERO; digit2<=ZERO; digit3<=SIX; end
      16'd6005: begin digit0<=FIVE; digit1<=ZERO; digit2<=ZERO; digit3<=SIX; end
      16'd6006: begin digit0<=SIX; digit1<=ZERO; digit2<=ZERO; digit3<=SIX; end
      16'd6007: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ZERO; digit3<=SIX; end
      16'd6008: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ZERO; digit3<=SIX; end
      16'd6009: begin digit0<=NINE; digit1<=ZERO; digit2<=ZERO; digit3<=SIX; end
      16'd6010: begin digit0<=ZERO; digit1<=ONE; digit2<=ZERO; digit3<=SIX; end
      16'd6011: begin digit0<=ONE; digit1<=ONE; digit2<=ZERO; digit3<=SIX; end
      16'd6012: begin digit0<=TWO; digit1<=ONE; digit2<=ZERO; digit3<=SIX; end
      16'd6013: begin digit0<=THREE; digit1<=ONE; digit2<=ZERO; digit3<=SIX; end
      16'd6014: begin digit0<=FOUR; digit1<=ONE; digit2<=ZERO; digit3<=SIX; end
      16'd6015: begin digit0<=FIVE; digit1<=ONE; digit2<=ZERO; digit3<=SIX; end
      16'd6016: begin digit0<=SIX; digit1<=ONE; digit2<=ZERO; digit3<=SIX; end
      16'd6017: begin digit0<=SEVEN; digit1<=ONE; digit2<=ZERO; digit3<=SIX; end
      16'd6018: begin digit0<=EIGHT; digit1<=ONE; digit2<=ZERO; digit3<=SIX; end
      16'd6019: begin digit0<=NINE; digit1<=ONE; digit2<=ZERO; digit3<=SIX; end
      16'd6020: begin digit0<=ZERO; digit1<=TWO; digit2<=ZERO; digit3<=SIX; end
      16'd6021: begin digit0<=ONE; digit1<=TWO; digit2<=ZERO; digit3<=SIX; end
      16'd6022: begin digit0<=TWO; digit1<=TWO; digit2<=ZERO; digit3<=SIX; end
      16'd6023: begin digit0<=THREE; digit1<=TWO; digit2<=ZERO; digit3<=SIX; end
      16'd6024: begin digit0<=FOUR; digit1<=TWO; digit2<=ZERO; digit3<=SIX; end
      16'd6025: begin digit0<=FIVE; digit1<=TWO; digit2<=ZERO; digit3<=SIX; end
      16'd6026: begin digit0<=SIX; digit1<=TWO; digit2<=ZERO; digit3<=SIX; end
      16'd6027: begin digit0<=SEVEN; digit1<=TWO; digit2<=ZERO; digit3<=SIX; end
      16'd6028: begin digit0<=EIGHT; digit1<=TWO; digit2<=ZERO; digit3<=SIX; end
      16'd6029: begin digit0<=NINE; digit1<=TWO; digit2<=ZERO; digit3<=SIX; end
      16'd6030: begin digit0<=ZERO; digit1<=THREE; digit2<=ZERO; digit3<=SIX; end
      16'd6031: begin digit0<=ONE; digit1<=THREE; digit2<=ZERO; digit3<=SIX; end
      16'd6032: begin digit0<=TWO; digit1<=THREE; digit2<=ZERO; digit3<=SIX; end
      16'd6033: begin digit0<=THREE; digit1<=THREE; digit2<=ZERO; digit3<=SIX; end
      16'd6034: begin digit0<=FOUR; digit1<=THREE; digit2<=ZERO; digit3<=SIX; end
      16'd6035: begin digit0<=FIVE; digit1<=THREE; digit2<=ZERO; digit3<=SIX; end
      16'd6036: begin digit0<=SIX; digit1<=THREE; digit2<=ZERO; digit3<=SIX; end
      16'd6037: begin digit0<=SEVEN; digit1<=THREE; digit2<=ZERO; digit3<=SIX; end
      16'd6038: begin digit0<=EIGHT; digit1<=THREE; digit2<=ZERO; digit3<=SIX; end
      16'd6039: begin digit0<=NINE; digit1<=THREE; digit2<=ZERO; digit3<=SIX; end
      16'd6040: begin digit0<=ZERO; digit1<=FOUR; digit2<=ZERO; digit3<=SIX; end
      16'd6041: begin digit0<=ONE; digit1<=FOUR; digit2<=ZERO; digit3<=SIX; end
      16'd6042: begin digit0<=TWO; digit1<=FOUR; digit2<=ZERO; digit3<=SIX; end
      16'd6043: begin digit0<=THREE; digit1<=FOUR; digit2<=ZERO; digit3<=SIX; end
      16'd6044: begin digit0<=FOUR; digit1<=FOUR; digit2<=ZERO; digit3<=SIX; end
      16'd6045: begin digit0<=FIVE; digit1<=FOUR; digit2<=ZERO; digit3<=SIX; end
      16'd6046: begin digit0<=SIX; digit1<=FOUR; digit2<=ZERO; digit3<=SIX; end
      16'd6047: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ZERO; digit3<=SIX; end
      16'd6048: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ZERO; digit3<=SIX; end
      16'd6049: begin digit0<=NINE; digit1<=FOUR; digit2<=ZERO; digit3<=SIX; end
      16'd6050: begin digit0<=ZERO; digit1<=FIVE; digit2<=ZERO; digit3<=SIX; end
      16'd6051: begin digit0<=ONE; digit1<=FIVE; digit2<=ZERO; digit3<=SIX; end
      16'd6052: begin digit0<=TWO; digit1<=FIVE; digit2<=ZERO; digit3<=SIX; end
      16'd6053: begin digit0<=THREE; digit1<=FIVE; digit2<=ZERO; digit3<=SIX; end
      16'd6054: begin digit0<=FOUR; digit1<=FIVE; digit2<=ZERO; digit3<=SIX; end
      16'd6055: begin digit0<=FIVE; digit1<=FIVE; digit2<=ZERO; digit3<=SIX; end
      16'd6056: begin digit0<=SIX; digit1<=FIVE; digit2<=ZERO; digit3<=SIX; end
      16'd6057: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ZERO; digit3<=SIX; end
      16'd6058: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ZERO; digit3<=SIX; end
      16'd6059: begin digit0<=NINE; digit1<=FIVE; digit2<=ZERO; digit3<=SIX; end
      16'd6060: begin digit0<=ZERO; digit1<=SIX; digit2<=ZERO; digit3<=SIX; end
      16'd6061: begin digit0<=ONE; digit1<=SIX; digit2<=ZERO; digit3<=SIX; end
      16'd6062: begin digit0<=TWO; digit1<=SIX; digit2<=ZERO; digit3<=SIX; end
      16'd6063: begin digit0<=THREE; digit1<=SIX; digit2<=ZERO; digit3<=SIX; end
      16'd6064: begin digit0<=FOUR; digit1<=SIX; digit2<=ZERO; digit3<=SIX; end
      16'd6065: begin digit0<=FIVE; digit1<=SIX; digit2<=ZERO; digit3<=SIX; end
      16'd6066: begin digit0<=SIX; digit1<=SIX; digit2<=ZERO; digit3<=SIX; end
      16'd6067: begin digit0<=SEVEN; digit1<=SIX; digit2<=ZERO; digit3<=SIX; end
      16'd6068: begin digit0<=EIGHT; digit1<=SIX; digit2<=ZERO; digit3<=SIX; end
      16'd6069: begin digit0<=NINE; digit1<=SIX; digit2<=ZERO; digit3<=SIX; end
      16'd6070: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ZERO; digit3<=SIX; end
      16'd6071: begin digit0<=ONE; digit1<=SEVEN; digit2<=ZERO; digit3<=SIX; end
      16'd6072: begin digit0<=TWO; digit1<=SEVEN; digit2<=ZERO; digit3<=SIX; end
      16'd6073: begin digit0<=THREE; digit1<=SEVEN; digit2<=ZERO; digit3<=SIX; end
      16'd6074: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ZERO; digit3<=SIX; end
      16'd6075: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ZERO; digit3<=SIX; end
      16'd6076: begin digit0<=SIX; digit1<=SEVEN; digit2<=ZERO; digit3<=SIX; end
      16'd6077: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ZERO; digit3<=SIX; end
      16'd6078: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ZERO; digit3<=SIX; end
      16'd6079: begin digit0<=NINE; digit1<=SEVEN; digit2<=ZERO; digit3<=SIX; end
      16'd6080: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ZERO; digit3<=SIX; end
      16'd6081: begin digit0<=ONE; digit1<=EIGHT; digit2<=ZERO; digit3<=SIX; end
      16'd6082: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ZERO; digit3<=SIX; end
      16'd6083: begin digit0<=THREE; digit1<=EIGHT; digit2<=ZERO; digit3<=SIX; end
      16'd6084: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ZERO; digit3<=SIX; end
      16'd6085: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ZERO; digit3<=SIX; end
      16'd6086: begin digit0<=SIX; digit1<=EIGHT; digit2<=ZERO; digit3<=SIX; end
      16'd6087: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ZERO; digit3<=SIX; end
      16'd6088: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ZERO; digit3<=SIX; end
      16'd6089: begin digit0<=NINE; digit1<=EIGHT; digit2<=ZERO; digit3<=SIX; end
      16'd6090: begin digit0<=ZERO; digit1<=NINE; digit2<=ZERO; digit3<=SIX; end
      16'd6091: begin digit0<=ONE; digit1<=NINE; digit2<=ZERO; digit3<=SIX; end
      16'd6092: begin digit0<=ZERO; digit1<=NINE; digit2<=ZERO; digit3<=SIX; end
      16'd6093: begin digit0<=THREE; digit1<=NINE; digit2<=ZERO; digit3<=SIX; end
      16'd6094: begin digit0<=FOUR; digit1<=NINE; digit2<=ZERO; digit3<=SIX; end
      16'd6095: begin digit0<=FIVE; digit1<=NINE; digit2<=ZERO; digit3<=SIX; end
      16'd6096: begin digit0<=SIX; digit1<=NINE; digit2<=ZERO; digit3<=SIX; end
      16'd6097: begin digit0<=SEVEN; digit1<=NINE; digit2<=ZERO; digit3<=SIX; end
      16'd6098: begin digit0<=EIGHT; digit1<=NINE; digit2<=ZERO; digit3<=SIX; end
      16'd6099: begin digit0<=NINE; digit1<=NINE; digit2<=ZERO; digit3<=SIX; end
	  16'd6100: begin digit0<=ZERO; digit1<=ZERO; digit2<=ONE; digit3<=SIX; end
      16'd6101: begin digit0<=ONE; digit1<=ZERO; digit2<=ONE; digit3<=SIX; end
      16'd6102: begin digit0<=TWO; digit1<=ZERO; digit2<=ONE; digit3<=SIX; end
      16'd6103: begin digit0<=THREE; digit1<=ZERO; digit2<=ONE; digit3<=SIX; end
      16'd6104: begin digit0<=FOUR; digit1<=ZERO; digit2<=ONE; digit3<=SIX; end
      16'd6105: begin digit0<=FIVE; digit1<=ZERO; digit2<=ONE; digit3<=SIX; end
      16'd6106: begin digit0<=SIX; digit1<=ZERO; digit2<=ONE; digit3<=SIX; end
      16'd6107: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ONE; digit3<=SIX; end
      16'd6108: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ONE; digit3<=SIX; end
      16'd6109: begin digit0<=NINE; digit1<=ZERO; digit2<=ONE; digit3<=SIX; end
      16'd6110: begin digit0<=ZERO; digit1<=ONE; digit2<=ONE; digit3<=SIX; end
      16'd6111: begin digit0<=ONE; digit1<=ONE; digit2<=ONE; digit3<=SIX; end
      16'd6112: begin digit0<=TWO; digit1<=ONE; digit2<=ONE; digit3<=SIX; end
      16'd6113: begin digit0<=THREE; digit1<=ONE; digit2<=ONE; digit3<=SIX; end
      16'd6114: begin digit0<=FOUR; digit1<=ONE; digit2<=ONE; digit3<=SIX; end
      16'd6115: begin digit0<=FIVE; digit1<=ONE; digit2<=ONE; digit3<=SIX; end
      16'd6116: begin digit0<=SIX; digit1<=ONE; digit2<=ONE; digit3<=SIX; end
      16'd6117: begin digit0<=SEVEN; digit1<=ONE; digit2<=ONE; digit3<=SIX; end
      16'd6118: begin digit0<=EIGHT; digit1<=ONE; digit2<=ONE; digit3<=SIX; end
      16'd6119: begin digit0<=NINE; digit1<=ONE; digit2<=ONE; digit3<=SIX; end
      16'd6120: begin digit0<=ZERO; digit1<=TWO; digit2<=ONE; digit3<=SIX; end
      16'd6121: begin digit0<=ONE; digit1<=TWO; digit2<=ONE; digit3<=SIX; end
      16'd6122: begin digit0<=TWO; digit1<=TWO; digit2<=ONE; digit3<=SIX; end
      16'd6123: begin digit0<=THREE; digit1<=TWO; digit2<=ONE; digit3<=SIX; end
      16'd6124: begin digit0<=FOUR; digit1<=TWO; digit2<=ONE; digit3<=SIX; end
      16'd6125: begin digit0<=FIVE; digit1<=TWO; digit2<=ONE; digit3<=SIX; end
      16'd6126: begin digit0<=SIX; digit1<=TWO; digit2<=ONE; digit3<=SIX; end
      16'd6127: begin digit0<=SEVEN; digit1<=TWO; digit2<=ONE; digit3<=SIX; end
      16'd6128: begin digit0<=EIGHT; digit1<=TWO; digit2<=ONE; digit3<=SIX; end
      16'd6129: begin digit0<=NINE; digit1<=TWO; digit2<=ONE; digit3<=SIX; end
      16'd6130: begin digit0<=ZERO; digit1<=THREE; digit2<=ONE; digit3<=SIX; end
      16'd6131: begin digit0<=ONE; digit1<=THREE; digit2<=ONE; digit3<=SIX; end
      16'd6132: begin digit0<=TWO; digit1<=THREE; digit2<=ONE; digit3<=SIX; end
      16'd6133: begin digit0<=THREE; digit1<=THREE; digit2<=ONE; digit3<=SIX; end
      16'd6134: begin digit0<=FOUR; digit1<=THREE; digit2<=ONE; digit3<=SIX; end
      16'd6135: begin digit0<=FIVE; digit1<=THREE; digit2<=ONE; digit3<=SIX; end
      16'd6136: begin digit0<=SIX; digit1<=THREE; digit2<=ONE; digit3<=SIX; end
      16'd6137: begin digit0<=SEVEN; digit1<=THREE; digit2<=ONE; digit3<=SIX; end
      16'd6138: begin digit0<=EIGHT; digit1<=THREE; digit2<=ONE; digit3<=SIX; end
      16'd6139: begin digit0<=NINE; digit1<=THREE; digit2<=ONE; digit3<=SIX; end
      16'd6140: begin digit0<=ZERO; digit1<=FOUR; digit2<=ONE; digit3<=SIX; end
      16'd6141: begin digit0<=ONE; digit1<=FOUR; digit2<=ONE; digit3<=SIX; end
      16'd6142: begin digit0<=TWO; digit1<=FOUR; digit2<=ONE; digit3<=SIX; end
      16'd6143: begin digit0<=THREE; digit1<=FOUR; digit2<=ONE; digit3<=SIX; end
      16'd6144: begin digit0<=FOUR; digit1<=FOUR; digit2<=ONE; digit3<=SIX; end
      16'd6145: begin digit0<=FIVE; digit1<=FOUR; digit2<=ONE; digit3<=SIX; end
      16'd6146: begin digit0<=SIX; digit1<=FOUR; digit2<=ONE; digit3<=SIX; end
      16'd6147: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ONE; digit3<=SIX; end
      16'd6148: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ONE; digit3<=SIX; end
      16'd6149: begin digit0<=NINE; digit1<=FOUR; digit2<=ONE; digit3<=SIX; end
      16'd6150: begin digit0<=ZERO; digit1<=FIVE; digit2<=ONE; digit3<=SIX; end
      16'd6151: begin digit0<=ONE; digit1<=FIVE; digit2<=ONE; digit3<=SIX; end
      16'd6152: begin digit0<=TWO; digit1<=FIVE; digit2<=ONE; digit3<=SIX; end
      16'd6153: begin digit0<=THREE; digit1<=FIVE; digit2<=ONE; digit3<=SIX; end
      16'd6154: begin digit0<=FOUR; digit1<=FIVE; digit2<=ONE; digit3<=SIX; end
      16'd6155: begin digit0<=FIVE; digit1<=FIVE; digit2<=ONE; digit3<=SIX; end
      16'd6156: begin digit0<=SIX; digit1<=FIVE; digit2<=ONE; digit3<=SIX; end
      16'd6157: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ONE; digit3<=SIX; end
      16'd6158: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ONE; digit3<=SIX; end
      16'd6159: begin digit0<=NINE; digit1<=FIVE; digit2<=ONE; digit3<=SIX; end
      16'd6160: begin digit0<=ZERO; digit1<=SIX; digit2<=ONE; digit3<=SIX; end
      16'd6161: begin digit0<=ONE; digit1<=SIX; digit2<=ONE; digit3<=SIX; end
      16'd6162: begin digit0<=TWO; digit1<=SIX; digit2<=ONE; digit3<=SIX; end
      16'd6163: begin digit0<=THREE; digit1<=SIX; digit2<=ONE; digit3<=SIX; end
      16'd6164: begin digit0<=FOUR; digit1<=SIX; digit2<=ONE; digit3<=SIX; end
      16'd6165: begin digit0<=FIVE; digit1<=SIX; digit2<=ONE; digit3<=SIX; end
      16'd6166: begin digit0<=SIX; digit1<=SIX; digit2<=ONE; digit3<=SIX; end
      16'd6167: begin digit0<=SEVEN; digit1<=SIX; digit2<=ONE; digit3<=SIX; end
      16'd6168: begin digit0<=EIGHT; digit1<=SIX; digit2<=ONE; digit3<=SIX; end
      16'd6169: begin digit0<=NINE; digit1<=SIX; digit2<=ONE; digit3<=SIX; end
      16'd6170: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ONE; digit3<=SIX; end
      16'd6171: begin digit0<=ONE; digit1<=SEVEN; digit2<=ONE; digit3<=SIX; end
      16'd6172: begin digit0<=TWO; digit1<=SEVEN; digit2<=ONE; digit3<=SIX; end
      16'd6173: begin digit0<=THREE; digit1<=SEVEN; digit2<=ONE; digit3<=SIX; end
      16'd6174: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ONE; digit3<=SIX; end
      16'd6175: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ONE; digit3<=SIX; end
      16'd6176: begin digit0<=SIX; digit1<=SEVEN; digit2<=ONE; digit3<=SIX; end
      16'd6177: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ONE; digit3<=SIX; end
      16'd6178: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ONE; digit3<=SIX; end
      16'd6179: begin digit0<=NINE; digit1<=SEVEN; digit2<=ONE; digit3<=SIX; end
      16'd6180: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=SIX; end
      16'd6181: begin digit0<=ONE; digit1<=EIGHT; digit2<=ONE; digit3<=SIX; end
      16'd6182: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=SIX; end
      16'd6183: begin digit0<=THREE; digit1<=EIGHT; digit2<=ONE; digit3<=SIX; end
      16'd6184: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ONE; digit3<=SIX; end
      16'd6185: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ONE; digit3<=SIX; end
      16'd6186: begin digit0<=SIX; digit1<=EIGHT; digit2<=ONE; digit3<=SIX; end
      16'd6187: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ONE; digit3<=SIX; end
      16'd6188: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ONE; digit3<=SIX; end
      16'd6189: begin digit0<=NINE; digit1<=EIGHT; digit2<=ONE; digit3<=SIX; end
      16'd6190: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=SIX; end
      16'd6191: begin digit0<=ONE; digit1<=NINE; digit2<=ONE; digit3<=SIX; end
      16'd6192: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=SIX; end
      16'd6193: begin digit0<=THREE; digit1<=NINE; digit2<=ONE; digit3<=SIX; end
      16'd6194: begin digit0<=FOUR; digit1<=NINE; digit2<=ONE; digit3<=SIX; end
      16'd6195: begin digit0<=FIVE; digit1<=NINE; digit2<=ONE; digit3<=SIX; end
      16'd6196: begin digit0<=SIX; digit1<=NINE; digit2<=ONE; digit3<=SIX; end
      16'd6197: begin digit0<=SEVEN; digit1<=NINE; digit2<=ONE; digit3<=SIX; end
      16'd6198: begin digit0<=EIGHT; digit1<=NINE; digit2<=ONE; digit3<=SIX; end
      16'd6199: begin digit0<=NINE; digit1<=NINE; digit2<=ONE; digit3<=SIX; end
	  16'd6200: begin digit0<=ZERO; digit1<=ZERO; digit2<=TWO; digit3<=SIX; end
      16'd6201: begin digit0<=ONE; digit1<=ZERO; digit2<=TWO; digit3<=SIX; end
      16'd6202: begin digit0<=TWO; digit1<=ZERO; digit2<=TWO; digit3<=SIX; end
      16'd6203: begin digit0<=THREE; digit1<=ZERO; digit2<=TWO; digit3<=SIX; end
      16'd6204: begin digit0<=FOUR; digit1<=ZERO; digit2<=TWO; digit3<=SIX; end
      16'd6205: begin digit0<=FIVE; digit1<=ZERO; digit2<=TWO; digit3<=SIX; end
      16'd6206: begin digit0<=SIX; digit1<=ZERO; digit2<=TWO; digit3<=SIX; end
      16'd6207: begin digit0<=SEVEN; digit1<=ZERO; digit2<=TWO; digit3<=SIX; end
      16'd6208: begin digit0<=EIGHT; digit1<=ZERO; digit2<=TWO; digit3<=SIX; end
      16'd6209: begin digit0<=NINE; digit1<=ZERO; digit2<=TWO; digit3<=SIX; end
      16'd6210: begin digit0<=ZERO; digit1<=ONE; digit2<=TWO; digit3<=SIX; end
      16'd6211: begin digit0<=ONE; digit1<=ONE; digit2<=TWO; digit3<=SIX; end
      16'd6212: begin digit0<=TWO; digit1<=ONE; digit2<=TWO; digit3<=SIX; end
      16'd6213: begin digit0<=THREE; digit1<=ONE; digit2<=TWO; digit3<=SIX; end
      16'd6214: begin digit0<=FOUR; digit1<=ONE; digit2<=TWO; digit3<=SIX; end
      16'd6215: begin digit0<=FIVE; digit1<=ONE; digit2<=TWO; digit3<=SIX; end
      16'd6216: begin digit0<=SIX; digit1<=ONE; digit2<=TWO; digit3<=SIX; end
      16'd6217: begin digit0<=SEVEN; digit1<=ONE; digit2<=TWO; digit3<=SIX; end
      16'd6218: begin digit0<=EIGHT; digit1<=ONE; digit2<=TWO; digit3<=SIX; end
      16'd6219: begin digit0<=NINE; digit1<=ONE; digit2<=TWO; digit3<=SIX; end
      16'd6220: begin digit0<=ZERO; digit1<=TWO; digit2<=TWO; digit3<=SIX; end
      16'd6221: begin digit0<=ONE; digit1<=TWO; digit2<=TWO; digit3<=SIX; end
      16'd6222: begin digit0<=TWO; digit1<=TWO; digit2<=TWO; digit3<=SIX; end
      16'd6223: begin digit0<=THREE; digit1<=TWO; digit2<=TWO; digit3<=SIX; end
      16'd6224: begin digit0<=FOUR; digit1<=TWO; digit2<=TWO; digit3<=SIX; end
      16'd6225: begin digit0<=FIVE; digit1<=TWO; digit2<=TWO; digit3<=SIX; end
      16'd6226: begin digit0<=SIX; digit1<=TWO; digit2<=TWO; digit3<=SIX; end
      16'd6227: begin digit0<=SEVEN; digit1<=TWO; digit2<=TWO; digit3<=SIX; end
      16'd6228: begin digit0<=EIGHT; digit1<=TWO; digit2<=TWO; digit3<=SIX; end
      16'd6229: begin digit0<=NINE; digit1<=TWO; digit2<=TWO; digit3<=SIX; end
      16'd6230: begin digit0<=ZERO; digit1<=THREE; digit2<=TWO; digit3<=SIX; end
      16'd6231: begin digit0<=ONE; digit1<=THREE; digit2<=TWO; digit3<=SIX; end
      16'd6232: begin digit0<=TWO; digit1<=THREE; digit2<=TWO; digit3<=SIX; end
      16'd6233: begin digit0<=THREE; digit1<=THREE; digit2<=TWO; digit3<=SIX; end
      16'd6234: begin digit0<=FOUR; digit1<=THREE; digit2<=TWO; digit3<=SIX; end
      16'd6235: begin digit0<=FIVE; digit1<=THREE; digit2<=TWO; digit3<=SIX; end
      16'd6236: begin digit0<=SIX; digit1<=THREE; digit2<=TWO; digit3<=SIX; end
      16'd6237: begin digit0<=SEVEN; digit1<=THREE; digit2<=TWO; digit3<=SIX; end
      16'd6238: begin digit0<=EIGHT; digit1<=THREE; digit2<=TWO; digit3<=SIX; end
      16'd6239: begin digit0<=NINE; digit1<=THREE; digit2<=TWO; digit3<=SIX; end
      16'd6240: begin digit0<=ZERO; digit1<=FOUR; digit2<=TWO; digit3<=SIX; end
      16'd6241: begin digit0<=ONE; digit1<=FOUR; digit2<=TWO; digit3<=SIX; end
      16'd6242: begin digit0<=TWO; digit1<=FOUR; digit2<=TWO; digit3<=SIX; end
      16'd6243: begin digit0<=THREE; digit1<=FOUR; digit2<=TWO; digit3<=SIX; end
      16'd6244: begin digit0<=FOUR; digit1<=FOUR; digit2<=TWO; digit3<=SIX; end
      16'd6245: begin digit0<=FIVE; digit1<=FOUR; digit2<=TWO; digit3<=SIX; end
      16'd6246: begin digit0<=SIX; digit1<=FOUR; digit2<=TWO; digit3<=SIX; end
      16'd6247: begin digit0<=SEVEN; digit1<=FOUR; digit2<=TWO; digit3<=SIX; end
      16'd6248: begin digit0<=EIGHT; digit1<=FOUR; digit2<=TWO; digit3<=SIX; end
      16'd6249: begin digit0<=NINE; digit1<=FOUR; digit2<=TWO; digit3<=SIX; end
      16'd6250: begin digit0<=ZERO; digit1<=FIVE; digit2<=TWO; digit3<=SIX; end
      16'd6251: begin digit0<=ONE; digit1<=FIVE; digit2<=TWO; digit3<=SIX; end
      16'd6252: begin digit0<=TWO; digit1<=FIVE; digit2<=TWO; digit3<=SIX; end
      16'd6253: begin digit0<=THREE; digit1<=FIVE; digit2<=TWO; digit3<=SIX; end
      16'd6254: begin digit0<=FOUR; digit1<=FIVE; digit2<=TWO; digit3<=SIX; end
      16'd6255: begin digit0<=FIVE; digit1<=FIVE; digit2<=TWO; digit3<=SIX; end
      16'd6256: begin digit0<=SIX; digit1<=FIVE; digit2<=TWO; digit3<=SIX; end
      16'd6257: begin digit0<=SEVEN; digit1<=FIVE; digit2<=TWO; digit3<=SIX; end
      16'd6258: begin digit0<=EIGHT; digit1<=FIVE; digit2<=TWO; digit3<=SIX; end
      16'd6259: begin digit0<=NINE; digit1<=FIVE; digit2<=TWO; digit3<=SIX; end
      16'd6260: begin digit0<=ZERO; digit1<=SIX; digit2<=TWO; digit3<=SIX; end
      16'd6261: begin digit0<=ONE; digit1<=SIX; digit2<=TWO; digit3<=SIX; end
      16'd6262: begin digit0<=TWO; digit1<=SIX; digit2<=TWO; digit3<=SIX; end
      16'd6263: begin digit0<=THREE; digit1<=SIX; digit2<=TWO; digit3<=SIX; end
      16'd6264: begin digit0<=FOUR; digit1<=SIX; digit2<=TWO; digit3<=SIX; end
      16'd6265: begin digit0<=FIVE; digit1<=SIX; digit2<=TWO; digit3<=SIX; end
      16'd6266: begin digit0<=SIX; digit1<=SIX; digit2<=TWO; digit3<=SIX; end
      16'd6267: begin digit0<=SEVEN; digit1<=SIX; digit2<=TWO; digit3<=SIX; end
      16'd6268: begin digit0<=EIGHT; digit1<=SIX; digit2<=TWO; digit3<=SIX; end
      16'd6269: begin digit0<=NINE; digit1<=SIX; digit2<=TWO; digit3<=SIX; end
      16'd6270: begin digit0<=ZERO; digit1<=SEVEN; digit2<=TWO; digit3<=SIX; end
      16'd6271: begin digit0<=ONE; digit1<=SEVEN; digit2<=TWO; digit3<=SIX; end
      16'd6272: begin digit0<=TWO; digit1<=SEVEN; digit2<=TWO; digit3<=SIX; end
      16'd6273: begin digit0<=THREE; digit1<=SEVEN; digit2<=TWO; digit3<=SIX; end
      16'd6274: begin digit0<=FOUR; digit1<=SEVEN; digit2<=TWO; digit3<=SIX; end
      16'd6275: begin digit0<=FIVE; digit1<=SEVEN; digit2<=TWO; digit3<=SIX; end
      16'd6276: begin digit0<=SIX; digit1<=SEVEN; digit2<=TWO; digit3<=SIX; end
      16'd6277: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=TWO; digit3<=SIX; end
      16'd6278: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=TWO; digit3<=SIX; end
      16'd6279: begin digit0<=NINE; digit1<=SEVEN; digit2<=TWO; digit3<=SIX; end
      16'd6280: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=SIX; end
      16'd6281: begin digit0<=ONE; digit1<=EIGHT; digit2<=TWO; digit3<=SIX; end
      16'd6282: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=SIX; end
      16'd6283: begin digit0<=THREE; digit1<=EIGHT; digit2<=TWO; digit3<=SIX; end
      16'd6284: begin digit0<=FOUR; digit1<=EIGHT; digit2<=TWO; digit3<=SIX; end
      16'd6285: begin digit0<=FIVE; digit1<=EIGHT; digit2<=TWO; digit3<=SIX; end
      16'd6286: begin digit0<=SIX; digit1<=EIGHT; digit2<=TWO; digit3<=SIX; end
      16'd6287: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=TWO; digit3<=SIX; end
      16'd6288: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=TWO; digit3<=SIX; end
      16'd6289: begin digit0<=NINE; digit1<=EIGHT; digit2<=TWO; digit3<=SIX; end
      16'd6290: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=SIX; end
      16'd6291: begin digit0<=ONE; digit1<=NINE; digit2<=TWO; digit3<=SIX; end
      16'd6292: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=SIX; end
      16'd6293: begin digit0<=THREE; digit1<=NINE; digit2<=TWO; digit3<=SIX; end
      16'd6294: begin digit0<=FOUR; digit1<=NINE; digit2<=TWO; digit3<=SIX; end
      16'd6295: begin digit0<=FIVE; digit1<=NINE; digit2<=TWO; digit3<=SIX; end
      16'd6296: begin digit0<=SIX; digit1<=NINE; digit2<=TWO; digit3<=SIX; end
      16'd6297: begin digit0<=SEVEN; digit1<=NINE; digit2<=TWO; digit3<=SIX; end
      16'd6298: begin digit0<=EIGHT; digit1<=NINE; digit2<=TWO; digit3<=SIX; end
      16'd6299: begin digit0<=NINE; digit1<=NINE; digit2<=TWO; digit3<=SIX; end
	  16'd6300: begin digit0<=ZERO; digit1<=ZERO; digit2<=THREE; digit3<=SIX; end
      16'd6301: begin digit0<=ONE; digit1<=ZERO; digit2<=THREE; digit3<=SIX; end
      16'd6302: begin digit0<=TWO; digit1<=ZERO; digit2<=THREE; digit3<=SIX; end
      16'd6303: begin digit0<=THREE; digit1<=ZERO; digit2<=THREE; digit3<=SIX; end
      16'd6304: begin digit0<=FOUR; digit1<=ZERO; digit2<=THREE; digit3<=SIX; end
      16'd6305: begin digit0<=FIVE; digit1<=ZERO; digit2<=THREE; digit3<=SIX; end
      16'd6306: begin digit0<=SIX; digit1<=ZERO; digit2<=THREE; digit3<=SIX; end
      16'd6307: begin digit0<=SEVEN; digit1<=ZERO; digit2<=THREE; digit3<=SIX; end
      16'd6308: begin digit0<=EIGHT; digit1<=ZERO; digit2<=THREE; digit3<=SIX; end
      16'd6309: begin digit0<=NINE; digit1<=ZERO; digit2<=THREE; digit3<=SIX; end
      16'd6310: begin digit0<=ZERO; digit1<=ONE; digit2<=THREE; digit3<=SIX; end
      16'd6311: begin digit0<=ONE; digit1<=ONE; digit2<=THREE; digit3<=SIX; end
      16'd6312: begin digit0<=TWO; digit1<=ONE; digit2<=THREE; digit3<=SIX; end
      16'd6313: begin digit0<=THREE; digit1<=ONE; digit2<=THREE; digit3<=SIX; end
      16'd6314: begin digit0<=FOUR; digit1<=ONE; digit2<=THREE; digit3<=SIX; end
      16'd6315: begin digit0<=FIVE; digit1<=ONE; digit2<=THREE; digit3<=SIX; end
      16'd6316: begin digit0<=SIX; digit1<=ONE; digit2<=THREE; digit3<=SIX; end
      16'd6317: begin digit0<=SEVEN; digit1<=ONE; digit2<=THREE; digit3<=SIX; end
      16'd6318: begin digit0<=EIGHT; digit1<=ONE; digit2<=THREE; digit3<=SIX; end
      16'd6319: begin digit0<=NINE; digit1<=ONE; digit2<=THREE; digit3<=SIX; end
      16'd6320: begin digit0<=ZERO; digit1<=TWO; digit2<=THREE; digit3<=SIX; end
      16'd6321: begin digit0<=ONE; digit1<=TWO; digit2<=THREE; digit3<=SIX; end
      16'd6322: begin digit0<=TWO; digit1<=TWO; digit2<=THREE; digit3<=SIX; end
      16'd6323: begin digit0<=THREE; digit1<=TWO; digit2<=THREE; digit3<=SIX; end
      16'd6324: begin digit0<=FOUR; digit1<=TWO; digit2<=THREE; digit3<=SIX; end
      16'd6325: begin digit0<=FIVE; digit1<=TWO; digit2<=THREE; digit3<=SIX; end
      16'd6326: begin digit0<=SIX; digit1<=TWO; digit2<=THREE; digit3<=SIX; end
      16'd6327: begin digit0<=SEVEN; digit1<=TWO; digit2<=THREE; digit3<=SIX; end
      16'd6328: begin digit0<=EIGHT; digit1<=TWO; digit2<=THREE; digit3<=SIX; end
      16'd6329: begin digit0<=NINE; digit1<=TWO; digit2<=THREE; digit3<=SIX; end
      16'd6330: begin digit0<=ZERO; digit1<=THREE; digit2<=THREE; digit3<=SIX; end
      16'd6331: begin digit0<=ONE; digit1<=THREE; digit2<=THREE; digit3<=SIX; end
      16'd6332: begin digit0<=TWO; digit1<=THREE; digit2<=THREE; digit3<=SIX; end
      16'd6333: begin digit0<=THREE; digit1<=THREE; digit2<=THREE; digit3<=SIX; end
      16'd6334: begin digit0<=FOUR; digit1<=THREE; digit2<=THREE; digit3<=SIX; end
      16'd6335: begin digit0<=FIVE; digit1<=THREE; digit2<=THREE; digit3<=SIX; end
      16'd6336: begin digit0<=SIX; digit1<=THREE; digit2<=THREE; digit3<=SIX; end
      16'd6337: begin digit0<=SEVEN; digit1<=THREE; digit2<=THREE; digit3<=SIX; end
      16'd6338: begin digit0<=EIGHT; digit1<=THREE; digit2<=THREE; digit3<=SIX; end
      16'd6339: begin digit0<=NINE; digit1<=THREE; digit2<=THREE; digit3<=SIX; end
      16'd6340: begin digit0<=ZERO; digit1<=FOUR; digit2<=THREE; digit3<=SIX; end
      16'd6341: begin digit0<=ONE; digit1<=FOUR; digit2<=THREE; digit3<=SIX; end
      16'd6342: begin digit0<=TWO; digit1<=FOUR; digit2<=THREE; digit3<=SIX; end
      16'd6343: begin digit0<=THREE; digit1<=FOUR; digit2<=THREE; digit3<=SIX; end
      16'd6344: begin digit0<=FOUR; digit1<=FOUR; digit2<=THREE; digit3<=SIX; end
      16'd6345: begin digit0<=FIVE; digit1<=FOUR; digit2<=THREE; digit3<=SIX; end
      16'd6346: begin digit0<=SIX; digit1<=FOUR; digit2<=THREE; digit3<=SIX; end
      16'd6347: begin digit0<=SEVEN; digit1<=FOUR; digit2<=THREE; digit3<=SIX; end
      16'd6348: begin digit0<=EIGHT; digit1<=FOUR; digit2<=THREE; digit3<=SIX; end
      16'd6349: begin digit0<=NINE; digit1<=FOUR; digit2<=THREE; digit3<=SIX; end
      16'd6350: begin digit0<=ZERO; digit1<=FIVE; digit2<=THREE; digit3<=SIX; end
      16'd6351: begin digit0<=ONE; digit1<=FIVE; digit2<=THREE; digit3<=SIX; end
      16'd6352: begin digit0<=TWO; digit1<=FIVE; digit2<=THREE; digit3<=SIX; end
      16'd6353: begin digit0<=THREE; digit1<=FIVE; digit2<=THREE; digit3<=SIX; end
      16'd6354: begin digit0<=FOUR; digit1<=FIVE; digit2<=THREE; digit3<=SIX; end
      16'd6355: begin digit0<=FIVE; digit1<=FIVE; digit2<=THREE; digit3<=SIX; end
      16'd6356: begin digit0<=SIX; digit1<=FIVE; digit2<=THREE; digit3<=SIX; end
      16'd6357: begin digit0<=SEVEN; digit1<=FIVE; digit2<=THREE; digit3<=SIX; end
      16'd6358: begin digit0<=EIGHT; digit1<=FIVE; digit2<=THREE; digit3<=SIX; end
      16'd6359: begin digit0<=NINE; digit1<=FIVE; digit2<=THREE; digit3<=SIX; end
      16'd6360: begin digit0<=ZERO; digit1<=SIX; digit2<=THREE; digit3<=SIX; end
      16'd6361: begin digit0<=ONE; digit1<=SIX; digit2<=THREE; digit3<=SIX; end
      16'd6362: begin digit0<=TWO; digit1<=SIX; digit2<=THREE; digit3<=SIX; end
      16'd6363: begin digit0<=THREE; digit1<=SIX; digit2<=THREE; digit3<=SIX; end
      16'd6364: begin digit0<=FOUR; digit1<=SIX; digit2<=THREE; digit3<=SIX; end
      16'd6365: begin digit0<=FIVE; digit1<=SIX; digit2<=THREE; digit3<=SIX; end
      16'd6366: begin digit0<=SIX; digit1<=SIX; digit2<=THREE; digit3<=SIX; end
      16'd6367: begin digit0<=SEVEN; digit1<=SIX; digit2<=THREE; digit3<=SIX; end
      16'd6368: begin digit0<=EIGHT; digit1<=SIX; digit2<=THREE; digit3<=SIX; end
      16'd6369: begin digit0<=NINE; digit1<=SIX; digit2<=THREE; digit3<=SIX; end
      16'd6370: begin digit0<=ZERO; digit1<=SEVEN; digit2<=THREE; digit3<=SIX; end
      16'd6371: begin digit0<=ONE; digit1<=SEVEN; digit2<=THREE; digit3<=SIX; end
      16'd6372: begin digit0<=TWO; digit1<=SEVEN; digit2<=THREE; digit3<=SIX; end
      16'd6373: begin digit0<=THREE; digit1<=SEVEN; digit2<=THREE; digit3<=SIX; end
      16'd6374: begin digit0<=FOUR; digit1<=SEVEN; digit2<=THREE; digit3<=SIX; end
      16'd6375: begin digit0<=FIVE; digit1<=SEVEN; digit2<=THREE; digit3<=SIX; end
      16'd6376: begin digit0<=SIX; digit1<=SEVEN; digit2<=THREE; digit3<=SIX; end
      16'd6377: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=THREE; digit3<=SIX; end
      16'd6378: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=THREE; digit3<=SIX; end
      16'd6379: begin digit0<=NINE; digit1<=SEVEN; digit2<=THREE; digit3<=SIX; end
      16'd6380: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=SIX; end
      16'd6381: begin digit0<=ONE; digit1<=EIGHT; digit2<=THREE; digit3<=SIX; end
      16'd6382: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=SIX; end
      16'd6383: begin digit0<=THREE; digit1<=EIGHT; digit2<=THREE; digit3<=SIX; end
      16'd6384: begin digit0<=FOUR; digit1<=EIGHT; digit2<=THREE; digit3<=SIX; end
      16'd6385: begin digit0<=FIVE; digit1<=EIGHT; digit2<=THREE; digit3<=SIX; end
      16'd6386: begin digit0<=SIX; digit1<=EIGHT; digit2<=THREE; digit3<=SIX; end
      16'd6387: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=THREE; digit3<=SIX; end
      16'd6388: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=THREE; digit3<=SIX; end
      16'd6389: begin digit0<=NINE; digit1<=EIGHT; digit2<=THREE; digit3<=SIX; end
      16'd6390: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=SIX; end
      16'd6391: begin digit0<=ONE; digit1<=NINE; digit2<=THREE; digit3<=SIX; end
      16'd6392: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=SIX; end
      16'd6393: begin digit0<=THREE; digit1<=NINE; digit2<=THREE; digit3<=SIX; end
      16'd6394: begin digit0<=FOUR; digit1<=NINE; digit2<=THREE; digit3<=SIX; end
      16'd6395: begin digit0<=FIVE; digit1<=NINE; digit2<=THREE; digit3<=SIX; end
      16'd6396: begin digit0<=SIX; digit1<=NINE; digit2<=THREE; digit3<=SIX; end
      16'd6397: begin digit0<=SEVEN; digit1<=NINE; digit2<=THREE; digit3<=SIX; end
      16'd6398: begin digit0<=EIGHT; digit1<=NINE; digit2<=THREE; digit3<=SIX; end
      16'd6399: begin digit0<=NINE; digit1<=NINE; digit2<=THREE; digit3<=SIX; end
	  16'd6400: begin digit0<=ZERO; digit1<=ZERO; digit2<=FOUR; digit3<=SIX; end
      16'd6401: begin digit0<=ONE; digit1<=ZERO; digit2<=FOUR; digit3<=SIX; end
      16'd6402: begin digit0<=TWO; digit1<=ZERO; digit2<=FOUR; digit3<=SIX; end
      16'd6403: begin digit0<=THREE; digit1<=ZERO; digit2<=FOUR; digit3<=SIX; end
      16'd6404: begin digit0<=FOUR; digit1<=ZERO; digit2<=FOUR; digit3<=SIX; end
      16'd6405: begin digit0<=FIVE; digit1<=ZERO; digit2<=FOUR; digit3<=SIX; end
      16'd6406: begin digit0<=SIX; digit1<=ZERO; digit2<=FOUR; digit3<=SIX; end
      16'd6407: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FOUR; digit3<=SIX; end
      16'd6408: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FOUR; digit3<=SIX; end
      16'd6409: begin digit0<=NINE; digit1<=ZERO; digit2<=FOUR; digit3<=SIX; end
      16'd6410: begin digit0<=ZERO; digit1<=ONE; digit2<=FOUR; digit3<=SIX; end
      16'd6411: begin digit0<=ONE; digit1<=ONE; digit2<=FOUR; digit3<=SIX; end
      16'd6412: begin digit0<=TWO; digit1<=ONE; digit2<=FOUR; digit3<=SIX; end
      16'd6413: begin digit0<=THREE; digit1<=ONE; digit2<=FOUR; digit3<=SIX; end
      16'd6414: begin digit0<=FOUR; digit1<=ONE; digit2<=FOUR; digit3<=SIX; end
      16'd6415: begin digit0<=FIVE; digit1<=ONE; digit2<=FOUR; digit3<=SIX; end
      16'd6416: begin digit0<=SIX; digit1<=ONE; digit2<=FOUR; digit3<=SIX; end
      16'd6417: begin digit0<=SEVEN; digit1<=ONE; digit2<=FOUR; digit3<=SIX; end
      16'd6418: begin digit0<=EIGHT; digit1<=ONE; digit2<=FOUR; digit3<=SIX; end
      16'd6419: begin digit0<=NINE; digit1<=ONE; digit2<=FOUR; digit3<=SIX; end
      16'd6420: begin digit0<=ZERO; digit1<=TWO; digit2<=FOUR; digit3<=SIX; end
      16'd6421: begin digit0<=ONE; digit1<=TWO; digit2<=FOUR; digit3<=SIX; end
      16'd6422: begin digit0<=TWO; digit1<=TWO; digit2<=FOUR; digit3<=SIX; end
      16'd6423: begin digit0<=THREE; digit1<=TWO; digit2<=FOUR; digit3<=SIX; end
      16'd6424: begin digit0<=FOUR; digit1<=TWO; digit2<=FOUR; digit3<=SIX; end
      16'd6425: begin digit0<=FIVE; digit1<=TWO; digit2<=FOUR; digit3<=SIX; end
      16'd6426: begin digit0<=SIX; digit1<=TWO; digit2<=FOUR; digit3<=SIX; end
      16'd6427: begin digit0<=SEVEN; digit1<=TWO; digit2<=FOUR; digit3<=SIX; end
      16'd6428: begin digit0<=EIGHT; digit1<=TWO; digit2<=FOUR; digit3<=SIX; end
      16'd6429: begin digit0<=NINE; digit1<=TWO; digit2<=FOUR; digit3<=SIX; end
      16'd6430: begin digit0<=ZERO; digit1<=THREE; digit2<=FOUR; digit3<=SIX; end
      16'd6431: begin digit0<=ONE; digit1<=THREE; digit2<=FOUR; digit3<=SIX; end
      16'd6432: begin digit0<=TWO; digit1<=THREE; digit2<=FOUR; digit3<=SIX; end
      16'd6433: begin digit0<=THREE; digit1<=THREE; digit2<=FOUR; digit3<=SIX; end
      16'd6434: begin digit0<=FOUR; digit1<=THREE; digit2<=FOUR; digit3<=SIX; end
      16'd6435: begin digit0<=FIVE; digit1<=THREE; digit2<=FOUR; digit3<=SIX; end
      16'd6436: begin digit0<=SIX; digit1<=THREE; digit2<=FOUR; digit3<=SIX; end
      16'd6437: begin digit0<=SEVEN; digit1<=THREE; digit2<=FOUR; digit3<=SIX; end
      16'd6438: begin digit0<=EIGHT; digit1<=THREE; digit2<=FOUR; digit3<=SIX; end
      16'd6439: begin digit0<=NINE; digit1<=THREE; digit2<=FOUR; digit3<=SIX; end
      16'd6440: begin digit0<=ZERO; digit1<=FOUR; digit2<=FOUR; digit3<=SIX; end
      16'd6441: begin digit0<=ONE; digit1<=FOUR; digit2<=FOUR; digit3<=SIX; end
      16'd6442: begin digit0<=TWO; digit1<=FOUR; digit2<=FOUR; digit3<=SIX; end
      16'd6443: begin digit0<=THREE; digit1<=FOUR; digit2<=FOUR; digit3<=SIX; end
      16'd6444: begin digit0<=FOUR; digit1<=FOUR; digit2<=FOUR; digit3<=SIX; end
      16'd6445: begin digit0<=FIVE; digit1<=FOUR; digit2<=FOUR; digit3<=SIX; end
      16'd6446: begin digit0<=SIX; digit1<=FOUR; digit2<=FOUR; digit3<=SIX; end
      16'd6447: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FOUR; digit3<=SIX; end
      16'd6448: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FOUR; digit3<=SIX; end
      16'd6449: begin digit0<=NINE; digit1<=FOUR; digit2<=FOUR; digit3<=SIX; end
      16'd6450: begin digit0<=ZERO; digit1<=FIVE; digit2<=FOUR; digit3<=SIX; end
      16'd6451: begin digit0<=ONE; digit1<=FIVE; digit2<=FOUR; digit3<=SIX; end
      16'd6452: begin digit0<=TWO; digit1<=FIVE; digit2<=FOUR; digit3<=SIX; end
      16'd6453: begin digit0<=THREE; digit1<=FIVE; digit2<=FOUR; digit3<=SIX; end
      16'd6454: begin digit0<=FOUR; digit1<=FIVE; digit2<=FOUR; digit3<=SIX; end
      16'd6455: begin digit0<=FIVE; digit1<=FIVE; digit2<=FOUR; digit3<=SIX; end
      16'd6456: begin digit0<=SIX; digit1<=FIVE; digit2<=FOUR; digit3<=SIX; end
      16'd6457: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FOUR; digit3<=SIX; end
      16'd6458: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FOUR; digit3<=SIX; end
      16'd6459: begin digit0<=NINE; digit1<=FIVE; digit2<=FOUR; digit3<=SIX; end
      16'd6460: begin digit0<=ZERO; digit1<=SIX; digit2<=FOUR; digit3<=SIX; end
      16'd6461: begin digit0<=ONE; digit1<=SIX; digit2<=FOUR; digit3<=SIX; end
      16'd6462: begin digit0<=TWO; digit1<=SIX; digit2<=FOUR; digit3<=SIX; end
      16'd6463: begin digit0<=THREE; digit1<=SIX; digit2<=FOUR; digit3<=SIX; end
      16'd6464: begin digit0<=FOUR; digit1<=SIX; digit2<=FOUR; digit3<=SIX; end
      16'd6465: begin digit0<=FIVE; digit1<=SIX; digit2<=FOUR; digit3<=SIX; end
      16'd6466: begin digit0<=SIX; digit1<=SIX; digit2<=FOUR; digit3<=SIX; end
      16'd6467: begin digit0<=SEVEN; digit1<=SIX; digit2<=FOUR; digit3<=SIX; end
      16'd6468: begin digit0<=EIGHT; digit1<=SIX; digit2<=FOUR; digit3<=SIX; end
      16'd6469: begin digit0<=NINE; digit1<=SIX; digit2<=FOUR; digit3<=SIX; end
      16'd6470: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FOUR; digit3<=SIX; end
      16'd6471: begin digit0<=ONE; digit1<=SEVEN; digit2<=FOUR; digit3<=SIX; end
      16'd6472: begin digit0<=TWO; digit1<=SEVEN; digit2<=FOUR; digit3<=SIX; end
      16'd6473: begin digit0<=THREE; digit1<=SEVEN; digit2<=FOUR; digit3<=SIX; end
      16'd6474: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FOUR; digit3<=SIX; end
      16'd6475: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FOUR; digit3<=SIX; end
      16'd6476: begin digit0<=SIX; digit1<=SEVEN; digit2<=FOUR; digit3<=SIX; end
      16'd6477: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FOUR; digit3<=SIX; end
      16'd6478: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FOUR; digit3<=SIX; end
      16'd6479: begin digit0<=NINE; digit1<=SEVEN; digit2<=FOUR; digit3<=SIX; end
      16'd6480: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=SIX; end
      16'd6481: begin digit0<=ONE; digit1<=EIGHT; digit2<=FOUR; digit3<=SIX; end
      16'd6482: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=SIX; end
      16'd6483: begin digit0<=THREE; digit1<=EIGHT; digit2<=FOUR; digit3<=SIX; end
      16'd6484: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FOUR; digit3<=SIX; end
      16'd6485: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FOUR; digit3<=SIX; end
      16'd6486: begin digit0<=SIX; digit1<=EIGHT; digit2<=FOUR; digit3<=SIX; end
      16'd6487: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FOUR; digit3<=SIX; end
      16'd6488: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FOUR; digit3<=SIX; end
      16'd6489: begin digit0<=NINE; digit1<=EIGHT; digit2<=FOUR; digit3<=SIX; end
      16'd6490: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=SIX; end
      16'd6491: begin digit0<=ONE; digit1<=NINE; digit2<=FOUR; digit3<=SIX; end
      16'd6492: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=SIX; end
      16'd6493: begin digit0<=THREE; digit1<=NINE; digit2<=FOUR; digit3<=SIX; end
      16'd6494: begin digit0<=FOUR; digit1<=NINE; digit2<=FOUR; digit3<=SIX; end
      16'd6495: begin digit0<=FIVE; digit1<=NINE; digit2<=FOUR; digit3<=SIX; end
      16'd6496: begin digit0<=SIX; digit1<=NINE; digit2<=FOUR; digit3<=SIX; end
      16'd6497: begin digit0<=SEVEN; digit1<=NINE; digit2<=FOUR; digit3<=SIX; end
      16'd6498: begin digit0<=EIGHT; digit1<=NINE; digit2<=FOUR; digit3<=SIX; end
      16'd6499: begin digit0<=NINE; digit1<=NINE; digit2<=FOUR; digit3<=SIX; end
	  16'd6500: begin digit0<=ZERO; digit1<=ZERO; digit2<=FIVE; digit3<=SIX; end
      16'd6501: begin digit0<=ONE; digit1<=ZERO; digit2<=FIVE; digit3<=SIX; end
      16'd6502: begin digit0<=TWO; digit1<=ZERO; digit2<=FIVE; digit3<=SIX; end
      16'd6503: begin digit0<=THREE; digit1<=ZERO; digit2<=FIVE; digit3<=SIX; end
      16'd6504: begin digit0<=FOUR; digit1<=ZERO; digit2<=FIVE; digit3<=SIX; end
      16'd6505: begin digit0<=FIVE; digit1<=ZERO; digit2<=FIVE; digit3<=SIX; end
      16'd6506: begin digit0<=SIX; digit1<=ZERO; digit2<=FIVE; digit3<=SIX; end
      16'd6507: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FIVE; digit3<=SIX; end
      16'd6508: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FIVE; digit3<=SIX; end
      16'd6509: begin digit0<=NINE; digit1<=ZERO; digit2<=FIVE; digit3<=SIX; end
      16'd6510: begin digit0<=ZERO; digit1<=ONE; digit2<=FIVE; digit3<=SIX; end
      16'd6511: begin digit0<=ONE; digit1<=ONE; digit2<=FIVE; digit3<=SIX; end
      16'd6512: begin digit0<=TWO; digit1<=ONE; digit2<=FIVE; digit3<=SIX; end
      16'd6513: begin digit0<=THREE; digit1<=ONE; digit2<=FIVE; digit3<=SIX; end
      16'd6514: begin digit0<=FOUR; digit1<=ONE; digit2<=FIVE; digit3<=SIX; end
      16'd6515: begin digit0<=FIVE; digit1<=ONE; digit2<=FIVE; digit3<=SIX; end
      16'd6516: begin digit0<=SIX; digit1<=ONE; digit2<=FIVE; digit3<=SIX; end
      16'd6517: begin digit0<=SEVEN; digit1<=ONE; digit2<=FIVE; digit3<=SIX; end
      16'd6518: begin digit0<=EIGHT; digit1<=ONE; digit2<=FIVE; digit3<=SIX; end
      16'd6519: begin digit0<=NINE; digit1<=ONE; digit2<=FIVE; digit3<=SIX; end
      16'd6520: begin digit0<=ZERO; digit1<=TWO; digit2<=FIVE; digit3<=SIX; end
      16'd6521: begin digit0<=ONE; digit1<=TWO; digit2<=FIVE; digit3<=SIX; end
      16'd6522: begin digit0<=TWO; digit1<=TWO; digit2<=FIVE; digit3<=SIX; end
      16'd6523: begin digit0<=THREE; digit1<=TWO; digit2<=FIVE; digit3<=SIX; end
      16'd6524: begin digit0<=FOUR; digit1<=TWO; digit2<=FIVE; digit3<=SIX; end
      16'd6525: begin digit0<=FIVE; digit1<=TWO; digit2<=FIVE; digit3<=SIX; end
      16'd6526: begin digit0<=SIX; digit1<=TWO; digit2<=FIVE; digit3<=SIX; end
      16'd6527: begin digit0<=SEVEN; digit1<=TWO; digit2<=FIVE; digit3<=SIX; end
      16'd6528: begin digit0<=EIGHT; digit1<=TWO; digit2<=FIVE; digit3<=SIX; end
      16'd6529: begin digit0<=NINE; digit1<=TWO; digit2<=FIVE; digit3<=SIX; end
      16'd6530: begin digit0<=ZERO; digit1<=THREE; digit2<=FIVE; digit3<=SIX; end
      16'd6531: begin digit0<=ONE; digit1<=THREE; digit2<=FIVE; digit3<=SIX; end
      16'd6532: begin digit0<=TWO; digit1<=THREE; digit2<=FIVE; digit3<=SIX; end
      16'd6533: begin digit0<=THREE; digit1<=THREE; digit2<=FIVE; digit3<=SIX; end
      16'd6534: begin digit0<=FOUR; digit1<=THREE; digit2<=FIVE; digit3<=SIX; end
      16'd6535: begin digit0<=FIVE; digit1<=THREE; digit2<=FIVE; digit3<=SIX; end
      16'd6536: begin digit0<=SIX; digit1<=THREE; digit2<=FIVE; digit3<=SIX; end
      16'd6537: begin digit0<=SEVEN; digit1<=THREE; digit2<=FIVE; digit3<=SIX; end
      16'd6538: begin digit0<=EIGHT; digit1<=THREE; digit2<=FIVE; digit3<=SIX; end
      16'd6539: begin digit0<=NINE; digit1<=THREE; digit2<=FIVE; digit3<=SIX; end
      16'd6540: begin digit0<=ZERO; digit1<=FOUR; digit2<=FIVE; digit3<=SIX; end
      16'd6541: begin digit0<=ONE; digit1<=FOUR; digit2<=FIVE; digit3<=SIX; end
      16'd6542: begin digit0<=TWO; digit1<=FOUR; digit2<=FIVE; digit3<=SIX; end
      16'd6543: begin digit0<=THREE; digit1<=FOUR; digit2<=FIVE; digit3<=SIX; end
      16'd6544: begin digit0<=FOUR; digit1<=FOUR; digit2<=FIVE; digit3<=SIX; end
      16'd6545: begin digit0<=FIVE; digit1<=FOUR; digit2<=FIVE; digit3<=SIX; end
      16'd6546: begin digit0<=SIX; digit1<=FOUR; digit2<=FIVE; digit3<=SIX; end
      16'd6547: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FIVE; digit3<=SIX; end
      16'd6548: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FIVE; digit3<=SIX; end
      16'd6549: begin digit0<=NINE; digit1<=FOUR; digit2<=FIVE; digit3<=SIX; end
      16'd6550: begin digit0<=ZERO; digit1<=FIVE; digit2<=FIVE; digit3<=SIX; end
      16'd6551: begin digit0<=ONE; digit1<=FIVE; digit2<=FIVE; digit3<=SIX; end
      16'd6552: begin digit0<=TWO; digit1<=FIVE; digit2<=FIVE; digit3<=SIX; end
      16'd6553: begin digit0<=THREE; digit1<=FIVE; digit2<=FIVE; digit3<=SIX; end
      16'd6554: begin digit0<=FOUR; digit1<=FIVE; digit2<=FIVE; digit3<=SIX; end
      16'd6555: begin digit0<=FIVE; digit1<=FIVE; digit2<=FIVE; digit3<=SIX; end
      16'd6556: begin digit0<=SIX; digit1<=FIVE; digit2<=FIVE; digit3<=SIX; end
      16'd6557: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FIVE; digit3<=SIX; end
      16'd6558: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FIVE; digit3<=SIX; end
      16'd6559: begin digit0<=NINE; digit1<=FIVE; digit2<=FIVE; digit3<=SIX; end
      16'd6560: begin digit0<=ZERO; digit1<=SIX; digit2<=FIVE; digit3<=SIX; end
      16'd6561: begin digit0<=ONE; digit1<=SIX; digit2<=FIVE; digit3<=SIX; end
      16'd6562: begin digit0<=TWO; digit1<=SIX; digit2<=FIVE; digit3<=SIX; end
      16'd6563: begin digit0<=THREE; digit1<=SIX; digit2<=FIVE; digit3<=SIX; end
      16'd6564: begin digit0<=FOUR; digit1<=SIX; digit2<=FIVE; digit3<=SIX; end
      16'd6565: begin digit0<=FIVE; digit1<=SIX; digit2<=FIVE; digit3<=SIX; end
      16'd6566: begin digit0<=SIX; digit1<=SIX; digit2<=FIVE; digit3<=SIX; end
      16'd6567: begin digit0<=SEVEN; digit1<=SIX; digit2<=FIVE; digit3<=SIX; end
      16'd6568: begin digit0<=EIGHT; digit1<=SIX; digit2<=FIVE; digit3<=SIX; end
      16'd6569: begin digit0<=NINE; digit1<=SIX; digit2<=FIVE; digit3<=SIX; end
      16'd6570: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FIVE; digit3<=SIX; end
      16'd6571: begin digit0<=ONE; digit1<=SEVEN; digit2<=FIVE; digit3<=SIX; end
      16'd6572: begin digit0<=TWO; digit1<=SEVEN; digit2<=FIVE; digit3<=SIX; end
      16'd6573: begin digit0<=THREE; digit1<=SEVEN; digit2<=FIVE; digit3<=SIX; end
      16'd6574: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FIVE; digit3<=SIX; end
      16'd6575: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FIVE; digit3<=SIX; end
      16'd6576: begin digit0<=SIX; digit1<=SEVEN; digit2<=FIVE; digit3<=SIX; end
      16'd6577: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FIVE; digit3<=SIX; end
      16'd6578: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FIVE; digit3<=SIX; end
      16'd6579: begin digit0<=NINE; digit1<=SEVEN; digit2<=FIVE; digit3<=SIX; end
      16'd6580: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=SIX; end
      16'd6581: begin digit0<=ONE; digit1<=EIGHT; digit2<=FIVE; digit3<=SIX; end
      16'd6582: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=SIX; end
      16'd6583: begin digit0<=THREE; digit1<=EIGHT; digit2<=FIVE; digit3<=SIX; end
      16'd6584: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FIVE; digit3<=SIX; end
      16'd6585: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FIVE; digit3<=SIX; end
      16'd6586: begin digit0<=SIX; digit1<=EIGHT; digit2<=FIVE; digit3<=SIX; end
      16'd6587: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FIVE; digit3<=SIX; end
      16'd6588: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FIVE; digit3<=SIX; end
      16'd6589: begin digit0<=NINE; digit1<=EIGHT; digit2<=FIVE; digit3<=SIX; end
      16'd6590: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=SIX; end
      16'd6591: begin digit0<=ONE; digit1<=NINE; digit2<=FIVE; digit3<=SIX; end
      16'd6592: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=SIX; end
      16'd6593: begin digit0<=THREE; digit1<=NINE; digit2<=FIVE; digit3<=SIX; end
      16'd6594: begin digit0<=FOUR; digit1<=NINE; digit2<=FIVE; digit3<=SIX; end
      16'd6595: begin digit0<=FIVE; digit1<=NINE; digit2<=FIVE; digit3<=SIX; end
      16'd6596: begin digit0<=SIX; digit1<=NINE; digit2<=FIVE; digit3<=SIX; end
      16'd6597: begin digit0<=SEVEN; digit1<=NINE; digit2<=FIVE; digit3<=SIX; end
      16'd6598: begin digit0<=EIGHT; digit1<=NINE; digit2<=FIVE; digit3<=SIX; end
      16'd6599: begin digit0<=NINE; digit1<=NINE; digit2<=FIVE; digit3<=SIX; end
	  16'd6600: begin digit0<=ZERO; digit1<=ZERO; digit2<=SIX; digit3<=SIX; end
      16'd6601: begin digit0<=ONE; digit1<=ZERO; digit2<=SIX; digit3<=SIX; end
      16'd6602: begin digit0<=TWO; digit1<=ZERO; digit2<=SIX; digit3<=SIX; end
      16'd6603: begin digit0<=THREE; digit1<=ZERO; digit2<=SIX; digit3<=SIX; end
      16'd6604: begin digit0<=FOUR; digit1<=ZERO; digit2<=SIX; digit3<=SIX; end
      16'd6605: begin digit0<=FIVE; digit1<=ZERO; digit2<=SIX; digit3<=SIX; end
      16'd6606: begin digit0<=SIX; digit1<=ZERO; digit2<=SIX; digit3<=SIX; end
      16'd6607: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SIX; digit3<=SIX; end
      16'd6608: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SIX; digit3<=SIX; end
      16'd6609: begin digit0<=NINE; digit1<=ZERO; digit2<=SIX; digit3<=SIX; end
      16'd6610: begin digit0<=ZERO; digit1<=ONE; digit2<=SIX; digit3<=SIX; end
      16'd6611: begin digit0<=ONE; digit1<=ONE; digit2<=SIX; digit3<=SIX; end
      16'd6612: begin digit0<=TWO; digit1<=ONE; digit2<=SIX; digit3<=SIX; end
      16'd6613: begin digit0<=THREE; digit1<=ONE; digit2<=SIX; digit3<=SIX; end
      16'd6614: begin digit0<=FOUR; digit1<=ONE; digit2<=SIX; digit3<=SIX; end
      16'd6615: begin digit0<=FIVE; digit1<=ONE; digit2<=SIX; digit3<=SIX; end
      16'd6616: begin digit0<=SIX; digit1<=ONE; digit2<=SIX; digit3<=SIX; end
      16'd6617: begin digit0<=SEVEN; digit1<=ONE; digit2<=SIX; digit3<=SIX; end
      16'd6618: begin digit0<=EIGHT; digit1<=ONE; digit2<=SIX; digit3<=SIX; end
      16'd6619: begin digit0<=NINE; digit1<=ONE; digit2<=SIX; digit3<=SIX; end
      16'd6620: begin digit0<=ZERO; digit1<=TWO; digit2<=SIX; digit3<=SIX; end
      16'd6621: begin digit0<=ONE; digit1<=TWO; digit2<=SIX; digit3<=SIX; end
      16'd6622: begin digit0<=TWO; digit1<=TWO; digit2<=SIX; digit3<=SIX; end
      16'd6623: begin digit0<=THREE; digit1<=TWO; digit2<=SIX; digit3<=SIX; end
      16'd6624: begin digit0<=FOUR; digit1<=TWO; digit2<=SIX; digit3<=SIX; end
      16'd6625: begin digit0<=FIVE; digit1<=TWO; digit2<=SIX; digit3<=SIX; end
      16'd6626: begin digit0<=SIX; digit1<=TWO; digit2<=SIX; digit3<=SIX; end
      16'd6627: begin digit0<=SEVEN; digit1<=TWO; digit2<=SIX; digit3<=SIX; end
      16'd6628: begin digit0<=EIGHT; digit1<=TWO; digit2<=SIX; digit3<=SIX; end
      16'd6629: begin digit0<=NINE; digit1<=TWO; digit2<=SIX; digit3<=SIX; end
      16'd6630: begin digit0<=ZERO; digit1<=THREE; digit2<=SIX; digit3<=SIX; end
      16'd6631: begin digit0<=ONE; digit1<=THREE; digit2<=SIX; digit3<=SIX; end
      16'd6632: begin digit0<=TWO; digit1<=THREE; digit2<=SIX; digit3<=SIX; end
      16'd6633: begin digit0<=THREE; digit1<=THREE; digit2<=SIX; digit3<=SIX; end
      16'd6634: begin digit0<=FOUR; digit1<=THREE; digit2<=SIX; digit3<=SIX; end
      16'd6635: begin digit0<=FIVE; digit1<=THREE; digit2<=SIX; digit3<=SIX; end
      16'd6636: begin digit0<=SIX; digit1<=THREE; digit2<=SIX; digit3<=SIX; end
      16'd6637: begin digit0<=SEVEN; digit1<=THREE; digit2<=SIX; digit3<=SIX; end
      16'd6638: begin digit0<=EIGHT; digit1<=THREE; digit2<=SIX; digit3<=SIX; end
      16'd6639: begin digit0<=NINE; digit1<=THREE; digit2<=SIX; digit3<=SIX; end
      16'd6640: begin digit0<=ZERO; digit1<=FOUR; digit2<=SIX; digit3<=SIX; end
      16'd6641: begin digit0<=ONE; digit1<=FOUR; digit2<=SIX; digit3<=SIX; end
      16'd6642: begin digit0<=TWO; digit1<=FOUR; digit2<=SIX; digit3<=SIX; end
      16'd6643: begin digit0<=THREE; digit1<=FOUR; digit2<=SIX; digit3<=SIX; end
      16'd6644: begin digit0<=FOUR; digit1<=FOUR; digit2<=SIX; digit3<=SIX; end
      16'd6645: begin digit0<=FIVE; digit1<=FOUR; digit2<=SIX; digit3<=SIX; end
      16'd6646: begin digit0<=SIX; digit1<=FOUR; digit2<=SIX; digit3<=SIX; end
      16'd6647: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SIX; digit3<=SIX; end
      16'd6648: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SIX; digit3<=SIX; end
      16'd6649: begin digit0<=NINE; digit1<=FOUR; digit2<=SIX; digit3<=SIX; end
      16'd6650: begin digit0<=ZERO; digit1<=FIVE; digit2<=SIX; digit3<=SIX; end
      16'd6651: begin digit0<=ONE; digit1<=FIVE; digit2<=SIX; digit3<=SIX; end
      16'd6652: begin digit0<=TWO; digit1<=FIVE; digit2<=SIX; digit3<=SIX; end
      16'd6653: begin digit0<=THREE; digit1<=FIVE; digit2<=SIX; digit3<=SIX; end
      16'd6654: begin digit0<=FOUR; digit1<=FIVE; digit2<=SIX; digit3<=SIX; end
      16'd6655: begin digit0<=FIVE; digit1<=FIVE; digit2<=SIX; digit3<=SIX; end
      16'd6656: begin digit0<=SIX; digit1<=FIVE; digit2<=SIX; digit3<=SIX; end
      16'd6657: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SIX; digit3<=SIX; end
      16'd6658: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SIX; digit3<=SIX; end
      16'd6659: begin digit0<=NINE; digit1<=FIVE; digit2<=SIX; digit3<=SIX; end
      16'd6660: begin digit0<=ZERO; digit1<=SIX; digit2<=SIX; digit3<=SIX; end
      16'd6661: begin digit0<=ONE; digit1<=SIX; digit2<=SIX; digit3<=SIX; end
      16'd6662: begin digit0<=TWO; digit1<=SIX; digit2<=SIX; digit3<=SIX; end
      16'd6663: begin digit0<=THREE; digit1<=SIX; digit2<=SIX; digit3<=SIX; end
      16'd6664: begin digit0<=FOUR; digit1<=SIX; digit2<=SIX; digit3<=SIX; end
      16'd6665: begin digit0<=FIVE; digit1<=SIX; digit2<=SIX; digit3<=SIX; end
      16'd6666: begin digit0<=SIX; digit1<=SIX; digit2<=SIX; digit3<=SIX; end
      16'd6667: begin digit0<=SEVEN; digit1<=SIX; digit2<=SIX; digit3<=SIX; end
      16'd6668: begin digit0<=EIGHT; digit1<=SIX; digit2<=SIX; digit3<=SIX; end
      16'd6669: begin digit0<=NINE; digit1<=SIX; digit2<=SIX; digit3<=SIX; end
      16'd6670: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SIX; digit3<=SIX; end
      16'd6671: begin digit0<=ONE; digit1<=SEVEN; digit2<=SIX; digit3<=SIX; end
      16'd6672: begin digit0<=TWO; digit1<=SEVEN; digit2<=SIX; digit3<=SIX; end
      16'd6673: begin digit0<=THREE; digit1<=SEVEN; digit2<=SIX; digit3<=SIX; end
      16'd6674: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SIX; digit3<=SIX; end
      16'd6675: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SIX; digit3<=SIX; end
      16'd6676: begin digit0<=SIX; digit1<=SEVEN; digit2<=SIX; digit3<=SIX; end
      16'd6677: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SIX; digit3<=SIX; end
      16'd6678: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SIX; digit3<=SIX; end
      16'd6679: begin digit0<=NINE; digit1<=SEVEN; digit2<=SIX; digit3<=SIX; end
      16'd6680: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=SIX; end
      16'd6681: begin digit0<=ONE; digit1<=EIGHT; digit2<=SIX; digit3<=SIX; end
      16'd6682: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=SIX; end
      16'd6683: begin digit0<=THREE; digit1<=EIGHT; digit2<=SIX; digit3<=SIX; end
      16'd6684: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SIX; digit3<=SIX; end
      16'd6685: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SIX; digit3<=SIX; end
      16'd6686: begin digit0<=SIX; digit1<=EIGHT; digit2<=SIX; digit3<=SIX; end
      16'd6687: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SIX; digit3<=SIX; end
      16'd6688: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SIX; digit3<=SIX; end
      16'd6689: begin digit0<=NINE; digit1<=EIGHT; digit2<=SIX; digit3<=SIX; end
      16'd6690: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=SIX; end
      16'd6691: begin digit0<=ONE; digit1<=NINE; digit2<=SIX; digit3<=SIX; end
      16'd6692: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=SIX; end
      16'd6693: begin digit0<=THREE; digit1<=NINE; digit2<=SIX; digit3<=SIX; end
      16'd6694: begin digit0<=FOUR; digit1<=NINE; digit2<=SIX; digit3<=SIX; end
      16'd6695: begin digit0<=FIVE; digit1<=NINE; digit2<=SIX; digit3<=SIX; end
      16'd6696: begin digit0<=SIX; digit1<=NINE; digit2<=SIX; digit3<=SIX; end
      16'd6697: begin digit0<=SEVEN; digit1<=NINE; digit2<=SIX; digit3<=SIX; end
      16'd6698: begin digit0<=EIGHT; digit1<=NINE; digit2<=SIX; digit3<=SIX; end
      16'd6699: begin digit0<=NINE; digit1<=NINE; digit2<=SIX; digit3<=SIX; end
	  16'd6700: begin digit0<=ZERO; digit1<=ZERO; digit2<=SEVEN; digit3<=SIX; end
      16'd6701: begin digit0<=ONE; digit1<=ZERO; digit2<=SEVEN; digit3<=SIX; end
      16'd6702: begin digit0<=TWO; digit1<=ZERO; digit2<=SEVEN; digit3<=SIX; end
      16'd6703: begin digit0<=THREE; digit1<=ZERO; digit2<=SEVEN; digit3<=SIX; end
      16'd6704: begin digit0<=FOUR; digit1<=ZERO; digit2<=SEVEN; digit3<=SIX; end
      16'd6705: begin digit0<=FIVE; digit1<=ZERO; digit2<=SEVEN; digit3<=SIX; end
      16'd6706: begin digit0<=SIX; digit1<=ZERO; digit2<=SEVEN; digit3<=SIX; end
      16'd6707: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SEVEN; digit3<=SIX; end
      16'd6708: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SEVEN; digit3<=SIX; end
      16'd6709: begin digit0<=NINE; digit1<=ZERO; digit2<=SEVEN; digit3<=SIX; end
      16'd6710: begin digit0<=ZERO; digit1<=ONE; digit2<=SEVEN; digit3<=SIX; end
      16'd6711: begin digit0<=ONE; digit1<=ONE; digit2<=SEVEN; digit3<=SIX; end
      16'd6712: begin digit0<=TWO; digit1<=ONE; digit2<=SEVEN; digit3<=SIX; end
      16'd6713: begin digit0<=THREE; digit1<=ONE; digit2<=SEVEN; digit3<=SIX; end
      16'd6714: begin digit0<=FOUR; digit1<=ONE; digit2<=SEVEN; digit3<=SIX; end
      16'd6715: begin digit0<=FIVE; digit1<=ONE; digit2<=SEVEN; digit3<=SIX; end
      16'd6716: begin digit0<=SIX; digit1<=ONE; digit2<=SEVEN; digit3<=SIX; end
      16'd6717: begin digit0<=SEVEN; digit1<=ONE; digit2<=SEVEN; digit3<=SIX; end
      16'd6718: begin digit0<=EIGHT; digit1<=ONE; digit2<=SEVEN; digit3<=SIX; end
      16'd6719: begin digit0<=NINE; digit1<=ONE; digit2<=SEVEN; digit3<=SIX; end
      16'd6720: begin digit0<=ZERO; digit1<=TWO; digit2<=SEVEN; digit3<=SIX; end
      16'd6721: begin digit0<=ONE; digit1<=TWO; digit2<=SEVEN; digit3<=SIX; end
      16'd6722: begin digit0<=TWO; digit1<=TWO; digit2<=SEVEN; digit3<=SIX; end
      16'd6723: begin digit0<=THREE; digit1<=TWO; digit2<=SEVEN; digit3<=SIX; end
      16'd6724: begin digit0<=FOUR; digit1<=TWO; digit2<=SEVEN; digit3<=SIX; end
      16'd6725: begin digit0<=FIVE; digit1<=TWO; digit2<=SEVEN; digit3<=SIX; end
      16'd6726: begin digit0<=SIX; digit1<=TWO; digit2<=SEVEN; digit3<=SIX; end
      16'd6727: begin digit0<=SEVEN; digit1<=TWO; digit2<=SEVEN; digit3<=SIX; end
      16'd6728: begin digit0<=EIGHT; digit1<=TWO; digit2<=SEVEN; digit3<=SIX; end
      16'd6729: begin digit0<=NINE; digit1<=TWO; digit2<=SEVEN; digit3<=SIX; end
      16'd6730: begin digit0<=ZERO; digit1<=THREE; digit2<=SEVEN; digit3<=SIX; end
      16'd6731: begin digit0<=ONE; digit1<=THREE; digit2<=SEVEN; digit3<=SIX; end
      16'd6732: begin digit0<=TWO; digit1<=THREE; digit2<=SEVEN; digit3<=SIX; end
      16'd6733: begin digit0<=THREE; digit1<=THREE; digit2<=SEVEN; digit3<=SIX; end
      16'd6734: begin digit0<=FOUR; digit1<=THREE; digit2<=SEVEN; digit3<=SIX; end
      16'd6735: begin digit0<=FIVE; digit1<=THREE; digit2<=SEVEN; digit3<=SIX; end
      16'd6736: begin digit0<=SIX; digit1<=THREE; digit2<=SEVEN; digit3<=SIX; end
      16'd6737: begin digit0<=SEVEN; digit1<=THREE; digit2<=SEVEN; digit3<=SIX; end
      16'd6738: begin digit0<=EIGHT; digit1<=THREE; digit2<=SEVEN; digit3<=SIX; end
      16'd6739: begin digit0<=NINE; digit1<=THREE; digit2<=SEVEN; digit3<=SIX; end
      16'd6740: begin digit0<=ZERO; digit1<=FOUR; digit2<=SEVEN; digit3<=SIX; end
      16'd6741: begin digit0<=ONE; digit1<=FOUR; digit2<=SEVEN; digit3<=SIX; end
      16'd6742: begin digit0<=TWO; digit1<=FOUR; digit2<=SEVEN; digit3<=SIX; end
      16'd6743: begin digit0<=THREE; digit1<=FOUR; digit2<=SEVEN; digit3<=SIX; end
      16'd6744: begin digit0<=FOUR; digit1<=FOUR; digit2<=SEVEN; digit3<=SIX; end
      16'd6745: begin digit0<=FIVE; digit1<=FOUR; digit2<=SEVEN; digit3<=SIX; end
      16'd6746: begin digit0<=SIX; digit1<=FOUR; digit2<=SEVEN; digit3<=SIX; end
      16'd6747: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SEVEN; digit3<=SIX; end
      16'd6748: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SEVEN; digit3<=SIX; end
      16'd6749: begin digit0<=NINE; digit1<=FOUR; digit2<=SEVEN; digit3<=SIX; end
      16'd6750: begin digit0<=ZERO; digit1<=FIVE; digit2<=SEVEN; digit3<=SIX; end
      16'd6751: begin digit0<=ONE; digit1<=FIVE; digit2<=SEVEN; digit3<=SIX; end
      16'd6752: begin digit0<=TWO; digit1<=FIVE; digit2<=SEVEN; digit3<=SIX; end
      16'd6753: begin digit0<=THREE; digit1<=FIVE; digit2<=SEVEN; digit3<=SIX; end
      16'd6754: begin digit0<=FOUR; digit1<=FIVE; digit2<=SEVEN; digit3<=SIX; end
      16'd6755: begin digit0<=FIVE; digit1<=FIVE; digit2<=SEVEN; digit3<=SIX; end
      16'd6756: begin digit0<=SIX; digit1<=FIVE; digit2<=SEVEN; digit3<=SIX; end
      16'd6757: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SEVEN; digit3<=SIX; end
      16'd6758: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SEVEN; digit3<=SIX; end
      16'd6759: begin digit0<=NINE; digit1<=FIVE; digit2<=SEVEN; digit3<=SIX; end
      16'd6760: begin digit0<=ZERO; digit1<=SIX; digit2<=SEVEN; digit3<=SIX; end
      16'd6761: begin digit0<=ONE; digit1<=SIX; digit2<=SEVEN; digit3<=SIX; end
      16'd6762: begin digit0<=TWO; digit1<=SIX; digit2<=SEVEN; digit3<=SIX; end
      16'd6763: begin digit0<=THREE; digit1<=SIX; digit2<=SEVEN; digit3<=SIX; end
      16'd6764: begin digit0<=FOUR; digit1<=SIX; digit2<=SEVEN; digit3<=SIX; end
      16'd6765: begin digit0<=FIVE; digit1<=SIX; digit2<=SEVEN; digit3<=SIX; end
      16'd6766: begin digit0<=SIX; digit1<=SIX; digit2<=SEVEN; digit3<=SIX; end
      16'd6767: begin digit0<=SEVEN; digit1<=SIX; digit2<=SEVEN; digit3<=SIX; end
      16'd6768: begin digit0<=EIGHT; digit1<=SIX; digit2<=SEVEN; digit3<=SIX; end
      16'd6769: begin digit0<=NINE; digit1<=SIX; digit2<=SEVEN; digit3<=SIX; end
      16'd6770: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SEVEN; digit3<=SIX; end
      16'd6771: begin digit0<=ONE; digit1<=SEVEN; digit2<=SEVEN; digit3<=SIX; end
      16'd6772: begin digit0<=TWO; digit1<=SEVEN; digit2<=SEVEN; digit3<=SIX; end
      16'd6773: begin digit0<=THREE; digit1<=SEVEN; digit2<=SEVEN; digit3<=SIX; end
      16'd6774: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SEVEN; digit3<=SIX; end
      16'd6775: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SEVEN; digit3<=SIX; end
      16'd6776: begin digit0<=SIX; digit1<=SEVEN; digit2<=SEVEN; digit3<=SIX; end
      16'd6777: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SEVEN; digit3<=SIX; end
      16'd6778: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SEVEN; digit3<=SIX; end
      16'd6779: begin digit0<=NINE; digit1<=SEVEN; digit2<=SEVEN; digit3<=SIX; end
      16'd6780: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=SIX; end
      16'd6781: begin digit0<=ONE; digit1<=EIGHT; digit2<=SEVEN; digit3<=SIX; end
      16'd6782: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=SIX; end
      16'd6783: begin digit0<=THREE; digit1<=EIGHT; digit2<=SEVEN; digit3<=SIX; end
      16'd6784: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SEVEN; digit3<=SIX; end
      16'd6785: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SEVEN; digit3<=SIX; end
      16'd6786: begin digit0<=SIX; digit1<=EIGHT; digit2<=SEVEN; digit3<=SIX; end
      16'd6787: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SEVEN; digit3<=SIX; end
      16'd6788: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SEVEN; digit3<=SIX; end
      16'd6789: begin digit0<=NINE; digit1<=EIGHT; digit2<=SEVEN; digit3<=SIX; end
      16'd6790: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=SIX; end
      16'd6791: begin digit0<=ONE; digit1<=NINE; digit2<=SEVEN; digit3<=SIX; end
      16'd6792: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=SIX; end
      16'd6793: begin digit0<=THREE; digit1<=NINE; digit2<=SEVEN; digit3<=SIX; end
      16'd6794: begin digit0<=FOUR; digit1<=NINE; digit2<=SEVEN; digit3<=SIX; end
      16'd6795: begin digit0<=FIVE; digit1<=NINE; digit2<=SEVEN; digit3<=SIX; end
      16'd6796: begin digit0<=SIX; digit1<=NINE; digit2<=SEVEN; digit3<=SIX; end
      16'd6797: begin digit0<=SEVEN; digit1<=NINE; digit2<=SEVEN; digit3<=SIX; end
      16'd6798: begin digit0<=EIGHT; digit1<=NINE; digit2<=SEVEN; digit3<=SIX; end
      16'd6799: begin digit0<=NINE; digit1<=NINE; digit2<=SEVEN; digit3<=SIX; end
	  16'd6800: begin digit0<=ZERO; digit1<=ZERO; digit2<=EIGHT; digit3<=SIX; end
      16'd6801: begin digit0<=ONE; digit1<=ZERO; digit2<=EIGHT; digit3<=SIX; end
      16'd6802: begin digit0<=TWO; digit1<=ZERO; digit2<=EIGHT; digit3<=SIX; end
      16'd6803: begin digit0<=THREE; digit1<=ZERO; digit2<=EIGHT; digit3<=SIX; end
      16'd6804: begin digit0<=FOUR; digit1<=ZERO; digit2<=EIGHT; digit3<=SIX; end
      16'd6805: begin digit0<=FIVE; digit1<=ZERO; digit2<=EIGHT; digit3<=SIX; end
      16'd6806: begin digit0<=SIX; digit1<=ZERO; digit2<=EIGHT; digit3<=SIX; end
      16'd6807: begin digit0<=SEVEN; digit1<=ZERO; digit2<=EIGHT; digit3<=SIX; end
      16'd6808: begin digit0<=EIGHT; digit1<=ZERO; digit2<=EIGHT; digit3<=SIX; end
      16'd6809: begin digit0<=NINE; digit1<=ZERO; digit2<=EIGHT; digit3<=SIX; end
      16'd6810: begin digit0<=ZERO; digit1<=ONE; digit2<=EIGHT; digit3<=SIX; end
      16'd6811: begin digit0<=ONE; digit1<=ONE; digit2<=EIGHT; digit3<=SIX; end
      16'd6812: begin digit0<=TWO; digit1<=ONE; digit2<=EIGHT; digit3<=SIX; end
      16'd6813: begin digit0<=THREE; digit1<=ONE; digit2<=EIGHT; digit3<=SIX; end
      16'd6814: begin digit0<=FOUR; digit1<=ONE; digit2<=EIGHT; digit3<=SIX; end
      16'd6815: begin digit0<=FIVE; digit1<=ONE; digit2<=EIGHT; digit3<=SIX; end
      16'd6816: begin digit0<=SIX; digit1<=ONE; digit2<=EIGHT; digit3<=SIX; end
      16'd6817: begin digit0<=SEVEN; digit1<=ONE; digit2<=EIGHT; digit3<=SIX; end
      16'd6818: begin digit0<=EIGHT; digit1<=ONE; digit2<=EIGHT; digit3<=SIX; end
      16'd6819: begin digit0<=NINE; digit1<=ONE; digit2<=EIGHT; digit3<=SIX; end
      16'd6820: begin digit0<=ZERO; digit1<=TWO; digit2<=EIGHT; digit3<=SIX; end
      16'd6821: begin digit0<=ONE; digit1<=TWO; digit2<=EIGHT; digit3<=SIX; end
      16'd6822: begin digit0<=TWO; digit1<=TWO; digit2<=EIGHT; digit3<=SIX; end
      16'd6823: begin digit0<=THREE; digit1<=TWO; digit2<=EIGHT; digit3<=SIX; end
      16'd6824: begin digit0<=FOUR; digit1<=TWO; digit2<=EIGHT; digit3<=SIX; end
      16'd6825: begin digit0<=FIVE; digit1<=TWO; digit2<=EIGHT; digit3<=SIX; end
      16'd6826: begin digit0<=SIX; digit1<=TWO; digit2<=EIGHT; digit3<=SIX; end
      16'd6827: begin digit0<=SEVEN; digit1<=TWO; digit2<=EIGHT; digit3<=SIX; end
      16'd6828: begin digit0<=EIGHT; digit1<=TWO; digit2<=EIGHT; digit3<=SIX; end
      16'd6829: begin digit0<=NINE; digit1<=TWO; digit2<=EIGHT; digit3<=SIX; end
      16'd6830: begin digit0<=ZERO; digit1<=THREE; digit2<=EIGHT; digit3<=SIX; end
      16'd6831: begin digit0<=ONE; digit1<=THREE; digit2<=EIGHT; digit3<=SIX; end
      16'd6832: begin digit0<=TWO; digit1<=THREE; digit2<=EIGHT; digit3<=SIX; end
      16'd6833: begin digit0<=THREE; digit1<=THREE; digit2<=EIGHT; digit3<=SIX; end
      16'd6834: begin digit0<=FOUR; digit1<=THREE; digit2<=EIGHT; digit3<=SIX; end
      16'd6835: begin digit0<=FIVE; digit1<=THREE; digit2<=EIGHT; digit3<=SIX; end
      16'd6836: begin digit0<=SIX; digit1<=THREE; digit2<=EIGHT; digit3<=SIX; end
      16'd6837: begin digit0<=SEVEN; digit1<=THREE; digit2<=EIGHT; digit3<=SIX; end
      16'd6838: begin digit0<=EIGHT; digit1<=THREE; digit2<=EIGHT; digit3<=SIX; end
      16'd6839: begin digit0<=NINE; digit1<=THREE; digit2<=EIGHT; digit3<=SIX; end
      16'd6840: begin digit0<=ZERO; digit1<=FOUR; digit2<=EIGHT; digit3<=SIX; end
      16'd6841: begin digit0<=ONE; digit1<=FOUR; digit2<=EIGHT; digit3<=SIX; end
      16'd6842: begin digit0<=TWO; digit1<=FOUR; digit2<=EIGHT; digit3<=SIX; end
      16'd6843: begin digit0<=THREE; digit1<=FOUR; digit2<=EIGHT; digit3<=SIX; end
      16'd6844: begin digit0<=FOUR; digit1<=FOUR; digit2<=EIGHT; digit3<=SIX; end
      16'd6845: begin digit0<=FIVE; digit1<=FOUR; digit2<=EIGHT; digit3<=SIX; end
      16'd6846: begin digit0<=SIX; digit1<=FOUR; digit2<=EIGHT; digit3<=SIX; end
      16'd6847: begin digit0<=SEVEN; digit1<=FOUR; digit2<=EIGHT; digit3<=SIX; end
      16'd6848: begin digit0<=EIGHT; digit1<=FOUR; digit2<=EIGHT; digit3<=SIX; end
      16'd6849: begin digit0<=NINE; digit1<=FOUR; digit2<=EIGHT; digit3<=SIX; end
      16'd6850: begin digit0<=ZERO; digit1<=FIVE; digit2<=EIGHT; digit3<=SIX; end
      16'd6851: begin digit0<=ONE; digit1<=FIVE; digit2<=EIGHT; digit3<=SIX; end
      16'd6852: begin digit0<=TWO; digit1<=FIVE; digit2<=EIGHT; digit3<=SIX; end
      16'd6853: begin digit0<=THREE; digit1<=FIVE; digit2<=EIGHT; digit3<=SIX; end
      16'd6854: begin digit0<=FOUR; digit1<=FIVE; digit2<=EIGHT; digit3<=SIX; end
      16'd6855: begin digit0<=FIVE; digit1<=FIVE; digit2<=EIGHT; digit3<=SIX; end
      16'd6856: begin digit0<=SIX; digit1<=FIVE; digit2<=EIGHT; digit3<=SIX; end
      16'd6857: begin digit0<=SEVEN; digit1<=FIVE; digit2<=EIGHT; digit3<=SIX; end
      16'd6858: begin digit0<=EIGHT; digit1<=FIVE; digit2<=EIGHT; digit3<=SIX; end
      16'd6859: begin digit0<=NINE; digit1<=FIVE; digit2<=EIGHT; digit3<=SIX; end
      16'd6860: begin digit0<=ZERO; digit1<=SIX; digit2<=EIGHT; digit3<=SIX; end
      16'd6861: begin digit0<=ONE; digit1<=SIX; digit2<=EIGHT; digit3<=SIX; end
      16'd6862: begin digit0<=TWO; digit1<=SIX; digit2<=EIGHT; digit3<=SIX; end
      16'd6863: begin digit0<=THREE; digit1<=SIX; digit2<=EIGHT; digit3<=SIX; end
      16'd6864: begin digit0<=FOUR; digit1<=SIX; digit2<=EIGHT; digit3<=SIX; end
      16'd6865: begin digit0<=FIVE; digit1<=SIX; digit2<=EIGHT; digit3<=SIX; end
      16'd6866: begin digit0<=SIX; digit1<=SIX; digit2<=EIGHT; digit3<=SIX; end
      16'd6867: begin digit0<=SEVEN; digit1<=SIX; digit2<=EIGHT; digit3<=SIX; end
      16'd6868: begin digit0<=EIGHT; digit1<=SIX; digit2<=EIGHT; digit3<=SIX; end
      16'd6869: begin digit0<=NINE; digit1<=SIX; digit2<=EIGHT; digit3<=SIX; end
      16'd6870: begin digit0<=ZERO; digit1<=SEVEN; digit2<=EIGHT; digit3<=SIX; end
      16'd6871: begin digit0<=ONE; digit1<=SEVEN; digit2<=EIGHT; digit3<=SIX; end
      16'd6872: begin digit0<=TWO; digit1<=SEVEN; digit2<=EIGHT; digit3<=SIX; end
      16'd6873: begin digit0<=THREE; digit1<=SEVEN; digit2<=EIGHT; digit3<=SIX; end
      16'd6874: begin digit0<=FOUR; digit1<=SEVEN; digit2<=EIGHT; digit3<=SIX; end
      16'd6875: begin digit0<=FIVE; digit1<=SEVEN; digit2<=EIGHT; digit3<=SIX; end
      16'd6876: begin digit0<=SIX; digit1<=SEVEN; digit2<=EIGHT; digit3<=SIX; end
      16'd6877: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=EIGHT; digit3<=SIX; end
      16'd6878: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=EIGHT; digit3<=SIX; end
      16'd6879: begin digit0<=NINE; digit1<=SEVEN; digit2<=EIGHT; digit3<=SIX; end
      16'd6880: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=SIX; end
      16'd6881: begin digit0<=ONE; digit1<=EIGHT; digit2<=EIGHT; digit3<=SIX; end
      16'd6882: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=SIX; end
      16'd6883: begin digit0<=THREE; digit1<=EIGHT; digit2<=EIGHT; digit3<=SIX; end
      16'd6884: begin digit0<=FOUR; digit1<=EIGHT; digit2<=EIGHT; digit3<=SIX; end
      16'd6885: begin digit0<=FIVE; digit1<=EIGHT; digit2<=EIGHT; digit3<=SIX; end
      16'd6886: begin digit0<=SIX; digit1<=EIGHT; digit2<=EIGHT; digit3<=SIX; end
      16'd6887: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=EIGHT; digit3<=SIX; end
      16'd6888: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=EIGHT; digit3<=SIX; end
      16'd6889: begin digit0<=NINE; digit1<=EIGHT; digit2<=EIGHT; digit3<=SIX; end
      16'd6890: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=SIX; end
      16'd6891: begin digit0<=ONE; digit1<=NINE; digit2<=EIGHT; digit3<=SIX; end
      16'd6892: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=SIX; end
      16'd6893: begin digit0<=THREE; digit1<=NINE; digit2<=EIGHT; digit3<=SIX; end
      16'd6894: begin digit0<=FOUR; digit1<=NINE; digit2<=EIGHT; digit3<=SIX; end
      16'd6895: begin digit0<=FIVE; digit1<=NINE; digit2<=EIGHT; digit3<=SIX; end
      16'd6896: begin digit0<=SIX; digit1<=NINE; digit2<=EIGHT; digit3<=SIX; end
      16'd6897: begin digit0<=SEVEN; digit1<=NINE; digit2<=EIGHT; digit3<=SIX; end
      16'd6898: begin digit0<=EIGHT; digit1<=NINE; digit2<=EIGHT; digit3<=SIX; end
      16'd6899: begin digit0<=NINE; digit1<=NINE; digit2<=EIGHT; digit3<=SIX; end
	  16'd6900: begin digit0<=ZERO; digit1<=ZERO; digit2<=NINE; digit3<=SIX; end
      16'd6901: begin digit0<=ONE; digit1<=ZERO; digit2<=NINE; digit3<=SIX; end
      16'd6902: begin digit0<=TWO; digit1<=ZERO; digit2<=NINE; digit3<=SIX; end
      16'd6903: begin digit0<=THREE; digit1<=ZERO; digit2<=NINE; digit3<=SIX; end
      16'd6904: begin digit0<=FOUR; digit1<=ZERO; digit2<=NINE; digit3<=SIX; end
      16'd6905: begin digit0<=FIVE; digit1<=ZERO; digit2<=NINE; digit3<=SIX; end
      16'd6906: begin digit0<=SIX; digit1<=ZERO; digit2<=NINE; digit3<=SIX; end
      16'd6907: begin digit0<=SEVEN; digit1<=ZERO; digit2<=NINE; digit3<=SIX; end
      16'd6908: begin digit0<=EIGHT; digit1<=ZERO; digit2<=NINE; digit3<=SIX; end
      16'd6909: begin digit0<=NINE; digit1<=ZERO; digit2<=NINE; digit3<=SIX; end
      16'd6910: begin digit0<=ZERO; digit1<=ONE; digit2<=NINE; digit3<=SIX; end
      16'd6911: begin digit0<=ONE; digit1<=ONE; digit2<=NINE; digit3<=SIX; end
      16'd6912: begin digit0<=TWO; digit1<=ONE; digit2<=NINE; digit3<=SIX; end
      16'd6913: begin digit0<=THREE; digit1<=ONE; digit2<=NINE; digit3<=SIX; end
      16'd6914: begin digit0<=FOUR; digit1<=ONE; digit2<=NINE; digit3<=SIX; end
      16'd6915: begin digit0<=FIVE; digit1<=ONE; digit2<=NINE; digit3<=SIX; end
      16'd6916: begin digit0<=SIX; digit1<=ONE; digit2<=NINE; digit3<=SIX; end
      16'd6917: begin digit0<=SEVEN; digit1<=ONE; digit2<=NINE; digit3<=SIX; end
      16'd6918: begin digit0<=EIGHT; digit1<=ONE; digit2<=NINE; digit3<=SIX; end
      16'd6919: begin digit0<=NINE; digit1<=ONE; digit2<=NINE; digit3<=SIX; end
      16'd6920: begin digit0<=ZERO; digit1<=TWO; digit2<=NINE; digit3<=SIX; end
      16'd6921: begin digit0<=ONE; digit1<=TWO; digit2<=NINE; digit3<=SIX; end
      16'd6922: begin digit0<=TWO; digit1<=TWO; digit2<=NINE; digit3<=SIX; end
      16'd6923: begin digit0<=THREE; digit1<=TWO; digit2<=NINE; digit3<=SIX; end
      16'd6924: begin digit0<=FOUR; digit1<=TWO; digit2<=NINE; digit3<=SIX; end
      16'd6925: begin digit0<=FIVE; digit1<=TWO; digit2<=NINE; digit3<=SIX; end
      16'd6926: begin digit0<=SIX; digit1<=TWO; digit2<=NINE; digit3<=SIX; end
      16'd6927: begin digit0<=SEVEN; digit1<=TWO; digit2<=NINE; digit3<=SIX; end
      16'd6928: begin digit0<=EIGHT; digit1<=TWO; digit2<=NINE; digit3<=SIX; end
      16'd6929: begin digit0<=NINE; digit1<=TWO; digit2<=NINE; digit3<=SIX; end
      16'd6930: begin digit0<=ZERO; digit1<=THREE; digit2<=NINE; digit3<=SIX; end
      16'd6931: begin digit0<=ONE; digit1<=THREE; digit2<=NINE; digit3<=SIX; end
      16'd6932: begin digit0<=TWO; digit1<=THREE; digit2<=NINE; digit3<=SIX; end
      16'd6933: begin digit0<=THREE; digit1<=THREE; digit2<=NINE; digit3<=SIX; end
      16'd6934: begin digit0<=FOUR; digit1<=THREE; digit2<=NINE; digit3<=SIX; end
      16'd6935: begin digit0<=FIVE; digit1<=THREE; digit2<=NINE; digit3<=SIX; end
      16'd6936: begin digit0<=SIX; digit1<=THREE; digit2<=NINE; digit3<=SIX; end
      16'd6937: begin digit0<=SEVEN; digit1<=THREE; digit2<=NINE; digit3<=SIX; end
      16'd6938: begin digit0<=EIGHT; digit1<=THREE; digit2<=NINE; digit3<=SIX; end
      16'd6939: begin digit0<=NINE; digit1<=THREE; digit2<=NINE; digit3<=SIX; end
      16'd6940: begin digit0<=ZERO; digit1<=FOUR; digit2<=NINE; digit3<=SIX; end
      16'd6941: begin digit0<=ONE; digit1<=FOUR; digit2<=NINE; digit3<=SIX; end
      16'd6942: begin digit0<=TWO; digit1<=FOUR; digit2<=NINE; digit3<=SIX; end
      16'd6943: begin digit0<=THREE; digit1<=FOUR; digit2<=NINE; digit3<=SIX; end
      16'd6944: begin digit0<=FOUR; digit1<=FOUR; digit2<=NINE; digit3<=SIX; end
      16'd6945: begin digit0<=FIVE; digit1<=FOUR; digit2<=NINE; digit3<=SIX; end
      16'd6946: begin digit0<=SIX; digit1<=FOUR; digit2<=NINE; digit3<=SIX; end
      16'd6947: begin digit0<=SEVEN; digit1<=FOUR; digit2<=NINE; digit3<=SIX; end
      16'd6948: begin digit0<=EIGHT; digit1<=FOUR; digit2<=NINE; digit3<=SIX; end
      16'd6949: begin digit0<=NINE; digit1<=FOUR; digit2<=NINE; digit3<=SIX; end
      16'd6950: begin digit0<=ZERO; digit1<=FIVE; digit2<=NINE; digit3<=SIX; end
      16'd6951: begin digit0<=ONE; digit1<=FIVE; digit2<=NINE; digit3<=SIX; end
      16'd6952: begin digit0<=TWO; digit1<=FIVE; digit2<=NINE; digit3<=SIX; end
      16'd6953: begin digit0<=THREE; digit1<=FIVE; digit2<=NINE; digit3<=SIX; end
      16'd6954: begin digit0<=FOUR; digit1<=FIVE; digit2<=NINE; digit3<=SIX; end
      16'd6955: begin digit0<=FIVE; digit1<=FIVE; digit2<=NINE; digit3<=SIX; end
      16'd6956: begin digit0<=SIX; digit1<=FIVE; digit2<=NINE; digit3<=SIX; end
      16'd6957: begin digit0<=SEVEN; digit1<=FIVE; digit2<=NINE; digit3<=SIX; end
      16'd6958: begin digit0<=EIGHT; digit1<=FIVE; digit2<=NINE; digit3<=SIX; end
      16'd6959: begin digit0<=NINE; digit1<=FIVE; digit2<=NINE; digit3<=SIX; end
      16'd6960: begin digit0<=ZERO; digit1<=SIX; digit2<=NINE; digit3<=SIX; end
      16'd6961: begin digit0<=ONE; digit1<=SIX; digit2<=NINE; digit3<=SIX; end
      16'd6962: begin digit0<=TWO; digit1<=SIX; digit2<=NINE; digit3<=SIX; end
      16'd6963: begin digit0<=THREE; digit1<=SIX; digit2<=NINE; digit3<=SIX; end
      16'd6964: begin digit0<=FOUR; digit1<=SIX; digit2<=NINE; digit3<=SIX; end
      16'd6965: begin digit0<=FIVE; digit1<=SIX; digit2<=NINE; digit3<=SIX; end
      16'd6966: begin digit0<=SIX; digit1<=SIX; digit2<=NINE; digit3<=SIX; end
      16'd6967: begin digit0<=SEVEN; digit1<=SIX; digit2<=NINE; digit3<=SIX; end
      16'd6968: begin digit0<=EIGHT; digit1<=SIX; digit2<=NINE; digit3<=SIX; end
      16'd6969: begin digit0<=NINE; digit1<=SIX; digit2<=NINE; digit3<=SIX; end
      16'd6970: begin digit0<=ZERO; digit1<=SEVEN; digit2<=NINE; digit3<=SIX; end
      16'd6971: begin digit0<=ONE; digit1<=SEVEN; digit2<=NINE; digit3<=SIX; end
      16'd6972: begin digit0<=TWO; digit1<=SEVEN; digit2<=NINE; digit3<=SIX; end
      16'd6973: begin digit0<=THREE; digit1<=SEVEN; digit2<=NINE; digit3<=SIX; end
      16'd6974: begin digit0<=FOUR; digit1<=SEVEN; digit2<=NINE; digit3<=SIX; end
      16'd6975: begin digit0<=FIVE; digit1<=SEVEN; digit2<=NINE; digit3<=SIX; end
      16'd6976: begin digit0<=SIX; digit1<=SEVEN; digit2<=NINE; digit3<=SIX; end
      16'd6977: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=NINE; digit3<=SIX; end
      16'd6978: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=NINE; digit3<=SIX; end
      16'd6979: begin digit0<=NINE; digit1<=SEVEN; digit2<=NINE; digit3<=SIX; end
      16'd6980: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=SIX; end
      16'd6981: begin digit0<=ONE; digit1<=EIGHT; digit2<=NINE; digit3<=SIX; end
      16'd6982: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=SIX; end
      16'd6983: begin digit0<=THREE; digit1<=EIGHT; digit2<=NINE; digit3<=SIX; end
      16'd6984: begin digit0<=FOUR; digit1<=EIGHT; digit2<=NINE; digit3<=SIX; end
      16'd6985: begin digit0<=FIVE; digit1<=EIGHT; digit2<=NINE; digit3<=SIX; end
      16'd6986: begin digit0<=SIX; digit1<=EIGHT; digit2<=NINE; digit3<=SIX; end
      16'd6987: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=NINE; digit3<=SIX; end
      16'd6988: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=NINE; digit3<=SIX; end
      16'd6989: begin digit0<=NINE; digit1<=EIGHT; digit2<=NINE; digit3<=SIX; end
      16'd6990: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=SIX; end
      16'd6991: begin digit0<=ONE; digit1<=NINE; digit2<=NINE; digit3<=SIX; end
      16'd6992: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=SIX; end
      16'd6993: begin digit0<=THREE; digit1<=NINE; digit2<=NINE; digit3<=SIX; end
      16'd6994: begin digit0<=FOUR; digit1<=NINE; digit2<=NINE; digit3<=SIX; end
      16'd6995: begin digit0<=FIVE; digit1<=NINE; digit2<=NINE; digit3<=SIX; end
      16'd6996: begin digit0<=SIX; digit1<=NINE; digit2<=NINE; digit3<=SIX; end
      16'd6997: begin digit0<=SEVEN; digit1<=NINE; digit2<=NINE; digit3<=SIX; end
      16'd6998: begin digit0<=EIGHT; digit1<=NINE; digit2<=NINE; digit3<=SIX; end
      16'd6999: begin digit0<=NINE; digit1<=NINE; digit2<=NINE; digit3<=SIX; end
	  16'd7000: begin digit0<=ZERO; digit1<=ZERO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7001: begin digit0<=ONE; digit1<=ZERO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7002: begin digit0<=TWO; digit1<=ZERO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7003: begin digit0<=THREE; digit1<=ZERO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7004: begin digit0<=FOUR; digit1<=ZERO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7005: begin digit0<=FIVE; digit1<=ZERO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7006: begin digit0<=SIX; digit1<=ZERO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7007: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7008: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7009: begin digit0<=NINE; digit1<=ZERO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7010: begin digit0<=ZERO; digit1<=ONE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7011: begin digit0<=ONE; digit1<=ONE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7012: begin digit0<=TWO; digit1<=ONE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7013: begin digit0<=THREE; digit1<=ONE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7014: begin digit0<=FOUR; digit1<=ONE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7015: begin digit0<=FIVE; digit1<=ONE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7016: begin digit0<=SIX; digit1<=ONE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7017: begin digit0<=SEVEN; digit1<=ONE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7018: begin digit0<=EIGHT; digit1<=ONE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7019: begin digit0<=NINE; digit1<=ONE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7020: begin digit0<=ZERO; digit1<=TWO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7021: begin digit0<=ONE; digit1<=TWO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7022: begin digit0<=TWO; digit1<=TWO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7023: begin digit0<=THREE; digit1<=TWO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7024: begin digit0<=FOUR; digit1<=TWO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7025: begin digit0<=FIVE; digit1<=TWO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7026: begin digit0<=SIX; digit1<=TWO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7027: begin digit0<=SEVEN; digit1<=TWO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7028: begin digit0<=EIGHT; digit1<=TWO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7029: begin digit0<=NINE; digit1<=TWO; digit2<=ZERO; digit3<=SEVEN; end
      16'd7030: begin digit0<=ZERO; digit1<=THREE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7031: begin digit0<=ONE; digit1<=THREE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7032: begin digit0<=TWO; digit1<=THREE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7033: begin digit0<=THREE; digit1<=THREE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7034: begin digit0<=FOUR; digit1<=THREE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7035: begin digit0<=FIVE; digit1<=THREE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7036: begin digit0<=SIX; digit1<=THREE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7037: begin digit0<=SEVEN; digit1<=THREE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7038: begin digit0<=EIGHT; digit1<=THREE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7039: begin digit0<=NINE; digit1<=THREE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7040: begin digit0<=ZERO; digit1<=FOUR; digit2<=ZERO; digit3<=SEVEN; end
      16'd7041: begin digit0<=ONE; digit1<=FOUR; digit2<=ZERO; digit3<=SEVEN; end
      16'd7042: begin digit0<=TWO; digit1<=FOUR; digit2<=ZERO; digit3<=SEVEN; end
      16'd7043: begin digit0<=THREE; digit1<=FOUR; digit2<=ZERO; digit3<=SEVEN; end
      16'd7044: begin digit0<=FOUR; digit1<=FOUR; digit2<=ZERO; digit3<=SEVEN; end
      16'd7045: begin digit0<=FIVE; digit1<=FOUR; digit2<=ZERO; digit3<=SEVEN; end
      16'd7046: begin digit0<=SIX; digit1<=FOUR; digit2<=ZERO; digit3<=SEVEN; end
      16'd7047: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ZERO; digit3<=SEVEN; end
      16'd7048: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ZERO; digit3<=SEVEN; end
      16'd7049: begin digit0<=NINE; digit1<=FOUR; digit2<=ZERO; digit3<=SEVEN; end
      16'd7050: begin digit0<=ZERO; digit1<=FIVE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7051: begin digit0<=ONE; digit1<=FIVE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7052: begin digit0<=TWO; digit1<=FIVE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7053: begin digit0<=THREE; digit1<=FIVE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7054: begin digit0<=FOUR; digit1<=FIVE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7055: begin digit0<=FIVE; digit1<=FIVE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7056: begin digit0<=SIX; digit1<=FIVE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7057: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7058: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7059: begin digit0<=NINE; digit1<=FIVE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7060: begin digit0<=ZERO; digit1<=SIX; digit2<=ZERO; digit3<=SEVEN; end
      16'd7061: begin digit0<=ONE; digit1<=SIX; digit2<=ZERO; digit3<=SEVEN; end
      16'd7062: begin digit0<=TWO; digit1<=SIX; digit2<=ZERO; digit3<=SEVEN; end
      16'd7063: begin digit0<=THREE; digit1<=SIX; digit2<=ZERO; digit3<=SEVEN; end
      16'd7064: begin digit0<=FOUR; digit1<=SIX; digit2<=ZERO; digit3<=SEVEN; end
      16'd7065: begin digit0<=FIVE; digit1<=SIX; digit2<=ZERO; digit3<=SEVEN; end
      16'd7066: begin digit0<=SIX; digit1<=SIX; digit2<=ZERO; digit3<=SEVEN; end
      16'd7067: begin digit0<=SEVEN; digit1<=SIX; digit2<=ZERO; digit3<=SEVEN; end
      16'd7068: begin digit0<=EIGHT; digit1<=SIX; digit2<=ZERO; digit3<=SEVEN; end
      16'd7069: begin digit0<=NINE; digit1<=SIX; digit2<=ZERO; digit3<=SEVEN; end
      16'd7070: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ZERO; digit3<=SEVEN; end
      16'd7071: begin digit0<=ONE; digit1<=SEVEN; digit2<=ZERO; digit3<=SEVEN; end
      16'd7072: begin digit0<=TWO; digit1<=SEVEN; digit2<=ZERO; digit3<=SEVEN; end
      16'd7073: begin digit0<=THREE; digit1<=SEVEN; digit2<=ZERO; digit3<=SEVEN; end
      16'd7074: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ZERO; digit3<=SEVEN; end
      16'd7075: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ZERO; digit3<=SEVEN; end
      16'd7076: begin digit0<=SIX; digit1<=SEVEN; digit2<=ZERO; digit3<=SEVEN; end
      16'd7077: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ZERO; digit3<=SEVEN; end
      16'd7078: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ZERO; digit3<=SEVEN; end
      16'd7079: begin digit0<=NINE; digit1<=SEVEN; digit2<=ZERO; digit3<=SEVEN; end
      16'd7080: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ZERO; digit3<=SEVEN; end
      16'd7081: begin digit0<=ONE; digit1<=EIGHT; digit2<=ZERO; digit3<=SEVEN; end
      16'd7082: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ZERO; digit3<=SEVEN; end
      16'd7083: begin digit0<=THREE; digit1<=EIGHT; digit2<=ZERO; digit3<=SEVEN; end
      16'd7084: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ZERO; digit3<=SEVEN; end
      16'd7085: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ZERO; digit3<=SEVEN; end
      16'd7086: begin digit0<=SIX; digit1<=EIGHT; digit2<=ZERO; digit3<=SEVEN; end
      16'd7087: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ZERO; digit3<=SEVEN; end
      16'd7088: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ZERO; digit3<=SEVEN; end
      16'd7089: begin digit0<=NINE; digit1<=EIGHT; digit2<=ZERO; digit3<=SEVEN; end
      16'd7090: begin digit0<=ZERO; digit1<=NINE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7091: begin digit0<=ONE; digit1<=NINE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7092: begin digit0<=ZERO; digit1<=NINE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7093: begin digit0<=THREE; digit1<=NINE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7094: begin digit0<=FOUR; digit1<=NINE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7095: begin digit0<=FIVE; digit1<=NINE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7096: begin digit0<=SIX; digit1<=NINE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7097: begin digit0<=SEVEN; digit1<=NINE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7098: begin digit0<=EIGHT; digit1<=NINE; digit2<=ZERO; digit3<=SEVEN; end
      16'd7099: begin digit0<=NINE; digit1<=NINE; digit2<=ZERO; digit3<=SEVEN; end
	  16'd7100: begin digit0<=ZERO; digit1<=ZERO; digit2<=ONE; digit3<=SEVEN; end
      16'd7101: begin digit0<=ONE; digit1<=ZERO; digit2<=ONE; digit3<=SEVEN; end
      16'd7102: begin digit0<=TWO; digit1<=ZERO; digit2<=ONE; digit3<=SEVEN; end
      16'd7103: begin digit0<=THREE; digit1<=ZERO; digit2<=ONE; digit3<=SEVEN; end
      16'd7104: begin digit0<=FOUR; digit1<=ZERO; digit2<=ONE; digit3<=SEVEN; end
      16'd7105: begin digit0<=FIVE; digit1<=ZERO; digit2<=ONE; digit3<=SEVEN; end
      16'd7106: begin digit0<=SIX; digit1<=ZERO; digit2<=ONE; digit3<=SEVEN; end
      16'd7107: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ONE; digit3<=SEVEN; end
      16'd7108: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ONE; digit3<=SEVEN; end
      16'd7109: begin digit0<=NINE; digit1<=ZERO; digit2<=ONE; digit3<=SEVEN; end
      16'd7110: begin digit0<=ZERO; digit1<=ONE; digit2<=ONE; digit3<=SEVEN; end
      16'd7111: begin digit0<=ONE; digit1<=ONE; digit2<=ONE; digit3<=SEVEN; end
      16'd7112: begin digit0<=TWO; digit1<=ONE; digit2<=ONE; digit3<=SEVEN; end
      16'd7113: begin digit0<=THREE; digit1<=ONE; digit2<=ONE; digit3<=SEVEN; end
      16'd7114: begin digit0<=FOUR; digit1<=ONE; digit2<=ONE; digit3<=SEVEN; end
      16'd7115: begin digit0<=FIVE; digit1<=ONE; digit2<=ONE; digit3<=SEVEN; end
      16'd7116: begin digit0<=SIX; digit1<=ONE; digit2<=ONE; digit3<=SEVEN; end
      16'd7117: begin digit0<=SEVEN; digit1<=ONE; digit2<=ONE; digit3<=SEVEN; end
      16'd7118: begin digit0<=EIGHT; digit1<=ONE; digit2<=ONE; digit3<=SEVEN; end
      16'd7119: begin digit0<=NINE; digit1<=ONE; digit2<=ONE; digit3<=SEVEN; end
      16'd7120: begin digit0<=ZERO; digit1<=TWO; digit2<=ONE; digit3<=SEVEN; end
      16'd7121: begin digit0<=ONE; digit1<=TWO; digit2<=ONE; digit3<=SEVEN; end
      16'd7122: begin digit0<=TWO; digit1<=TWO; digit2<=ONE; digit3<=SEVEN; end
      16'd7123: begin digit0<=THREE; digit1<=TWO; digit2<=ONE; digit3<=SEVEN; end
      16'd7124: begin digit0<=FOUR; digit1<=TWO; digit2<=ONE; digit3<=SEVEN; end
      16'd7125: begin digit0<=FIVE; digit1<=TWO; digit2<=ONE; digit3<=SEVEN; end
      16'd7126: begin digit0<=SIX; digit1<=TWO; digit2<=ONE; digit3<=SEVEN; end
      16'd7127: begin digit0<=SEVEN; digit1<=TWO; digit2<=ONE; digit3<=SEVEN; end
      16'd7128: begin digit0<=EIGHT; digit1<=TWO; digit2<=ONE; digit3<=SEVEN; end
      16'd7129: begin digit0<=NINE; digit1<=TWO; digit2<=ONE; digit3<=SEVEN; end
      16'd7130: begin digit0<=ZERO; digit1<=THREE; digit2<=ONE; digit3<=SEVEN; end
      16'd7131: begin digit0<=ONE; digit1<=THREE; digit2<=ONE; digit3<=SEVEN; end
      16'd7132: begin digit0<=TWO; digit1<=THREE; digit2<=ONE; digit3<=SEVEN; end
      16'd7133: begin digit0<=THREE; digit1<=THREE; digit2<=ONE; digit3<=SEVEN; end
      16'd7134: begin digit0<=FOUR; digit1<=THREE; digit2<=ONE; digit3<=SEVEN; end
      16'd7135: begin digit0<=FIVE; digit1<=THREE; digit2<=ONE; digit3<=SEVEN; end
      16'd7136: begin digit0<=SIX; digit1<=THREE; digit2<=ONE; digit3<=SEVEN; end
      16'd7137: begin digit0<=SEVEN; digit1<=THREE; digit2<=ONE; digit3<=SEVEN; end
      16'd7138: begin digit0<=EIGHT; digit1<=THREE; digit2<=ONE; digit3<=SEVEN; end
      16'd7139: begin digit0<=NINE; digit1<=THREE; digit2<=ONE; digit3<=SEVEN; end
      16'd7140: begin digit0<=ZERO; digit1<=FOUR; digit2<=ONE; digit3<=SEVEN; end
      16'd7141: begin digit0<=ONE; digit1<=FOUR; digit2<=ONE; digit3<=SEVEN; end
      16'd7142: begin digit0<=TWO; digit1<=FOUR; digit2<=ONE; digit3<=SEVEN; end
      16'd7143: begin digit0<=THREE; digit1<=FOUR; digit2<=ONE; digit3<=SEVEN; end
      16'd7144: begin digit0<=FOUR; digit1<=FOUR; digit2<=ONE; digit3<=SEVEN; end
      16'd7145: begin digit0<=FIVE; digit1<=FOUR; digit2<=ONE; digit3<=SEVEN; end
      16'd7146: begin digit0<=SIX; digit1<=FOUR; digit2<=ONE; digit3<=SEVEN; end
      16'd7147: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ONE; digit3<=SEVEN; end
      16'd7148: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ONE; digit3<=SEVEN; end
      16'd7149: begin digit0<=NINE; digit1<=FOUR; digit2<=ONE; digit3<=SEVEN; end
      16'd7150: begin digit0<=ZERO; digit1<=FIVE; digit2<=ONE; digit3<=SEVEN; end
      16'd7151: begin digit0<=ONE; digit1<=FIVE; digit2<=ONE; digit3<=SEVEN; end
      16'd7152: begin digit0<=TWO; digit1<=FIVE; digit2<=ONE; digit3<=SEVEN; end
      16'd7153: begin digit0<=THREE; digit1<=FIVE; digit2<=ONE; digit3<=SEVEN; end
      16'd7154: begin digit0<=FOUR; digit1<=FIVE; digit2<=ONE; digit3<=SEVEN; end
      16'd7155: begin digit0<=FIVE; digit1<=FIVE; digit2<=ONE; digit3<=SEVEN; end
      16'd7156: begin digit0<=SIX; digit1<=FIVE; digit2<=ONE; digit3<=SEVEN; end
      16'd7157: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ONE; digit3<=SEVEN; end
      16'd7158: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ONE; digit3<=SEVEN; end
      16'd7159: begin digit0<=NINE; digit1<=FIVE; digit2<=ONE; digit3<=SEVEN; end
      16'd7160: begin digit0<=ZERO; digit1<=SIX; digit2<=ONE; digit3<=SEVEN; end
      16'd7161: begin digit0<=ONE; digit1<=SIX; digit2<=ONE; digit3<=SEVEN; end
      16'd7162: begin digit0<=TWO; digit1<=SIX; digit2<=ONE; digit3<=SEVEN; end
      16'd7163: begin digit0<=THREE; digit1<=SIX; digit2<=ONE; digit3<=SEVEN; end
      16'd7164: begin digit0<=FOUR; digit1<=SIX; digit2<=ONE; digit3<=SEVEN; end
      16'd7165: begin digit0<=FIVE; digit1<=SIX; digit2<=ONE; digit3<=SEVEN; end
      16'd7166: begin digit0<=SIX; digit1<=SIX; digit2<=ONE; digit3<=SEVEN; end
      16'd7167: begin digit0<=SEVEN; digit1<=SIX; digit2<=ONE; digit3<=SEVEN; end
      16'd7168: begin digit0<=EIGHT; digit1<=SIX; digit2<=ONE; digit3<=SEVEN; end
      16'd7169: begin digit0<=NINE; digit1<=SIX; digit2<=ONE; digit3<=SEVEN; end
      16'd7170: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ONE; digit3<=SEVEN; end
      16'd7171: begin digit0<=ONE; digit1<=SEVEN; digit2<=ONE; digit3<=SEVEN; end
      16'd7172: begin digit0<=TWO; digit1<=SEVEN; digit2<=ONE; digit3<=SEVEN; end
      16'd7173: begin digit0<=THREE; digit1<=SEVEN; digit2<=ONE; digit3<=SEVEN; end
      16'd7174: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ONE; digit3<=SEVEN; end
      16'd7175: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ONE; digit3<=SEVEN; end
      16'd7176: begin digit0<=SIX; digit1<=SEVEN; digit2<=ONE; digit3<=SEVEN; end
      16'd7177: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ONE; digit3<=SEVEN; end
      16'd7178: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ONE; digit3<=SEVEN; end
      16'd7179: begin digit0<=NINE; digit1<=SEVEN; digit2<=ONE; digit3<=SEVEN; end
      16'd7180: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=SEVEN; end
      16'd7181: begin digit0<=ONE; digit1<=EIGHT; digit2<=ONE; digit3<=SEVEN; end
      16'd7182: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=SEVEN; end
      16'd7183: begin digit0<=THREE; digit1<=EIGHT; digit2<=ONE; digit3<=SEVEN; end
      16'd7184: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ONE; digit3<=SEVEN; end
      16'd7185: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ONE; digit3<=SEVEN; end
      16'd7186: begin digit0<=SIX; digit1<=EIGHT; digit2<=ONE; digit3<=SEVEN; end
      16'd7187: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ONE; digit3<=SEVEN; end
      16'd7188: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ONE; digit3<=SEVEN; end
      16'd7189: begin digit0<=NINE; digit1<=EIGHT; digit2<=ONE; digit3<=SEVEN; end
      16'd7190: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=SEVEN; end
      16'd7191: begin digit0<=ONE; digit1<=NINE; digit2<=ONE; digit3<=SEVEN; end
      16'd7192: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=SEVEN; end
      16'd7193: begin digit0<=THREE; digit1<=NINE; digit2<=ONE; digit3<=SEVEN; end
      16'd7194: begin digit0<=FOUR; digit1<=NINE; digit2<=ONE; digit3<=SEVEN; end
      16'd7195: begin digit0<=FIVE; digit1<=NINE; digit2<=ONE; digit3<=SEVEN; end
      16'd7196: begin digit0<=SIX; digit1<=NINE; digit2<=ONE; digit3<=SEVEN; end
      16'd7197: begin digit0<=SEVEN; digit1<=NINE; digit2<=ONE; digit3<=SEVEN; end
      16'd7198: begin digit0<=EIGHT; digit1<=NINE; digit2<=ONE; digit3<=SEVEN; end
      16'd7199: begin digit0<=NINE; digit1<=NINE; digit2<=ONE; digit3<=SEVEN; end
	  16'd7200: begin digit0<=ZERO; digit1<=ZERO; digit2<=TWO; digit3<=SEVEN; end
      16'd7201: begin digit0<=ONE; digit1<=ZERO; digit2<=TWO; digit3<=SEVEN; end
      16'd7202: begin digit0<=TWO; digit1<=ZERO; digit2<=TWO; digit3<=SEVEN; end
      16'd7203: begin digit0<=THREE; digit1<=ZERO; digit2<=TWO; digit3<=SEVEN; end
      16'd7204: begin digit0<=FOUR; digit1<=ZERO; digit2<=TWO; digit3<=SEVEN; end
      16'd7205: begin digit0<=FIVE; digit1<=ZERO; digit2<=TWO; digit3<=SEVEN; end
      16'd7206: begin digit0<=SIX; digit1<=ZERO; digit2<=TWO; digit3<=SEVEN; end
      16'd7207: begin digit0<=SEVEN; digit1<=ZERO; digit2<=TWO; digit3<=SEVEN; end
      16'd7208: begin digit0<=EIGHT; digit1<=ZERO; digit2<=TWO; digit3<=SEVEN; end
      16'd7209: begin digit0<=NINE; digit1<=ZERO; digit2<=TWO; digit3<=SEVEN; end
      16'd7210: begin digit0<=ZERO; digit1<=ONE; digit2<=TWO; digit3<=SEVEN; end
      16'd7211: begin digit0<=ONE; digit1<=ONE; digit2<=TWO; digit3<=SEVEN; end
      16'd7212: begin digit0<=TWO; digit1<=ONE; digit2<=TWO; digit3<=SEVEN; end
      16'd7213: begin digit0<=THREE; digit1<=ONE; digit2<=TWO; digit3<=SEVEN; end
      16'd7214: begin digit0<=FOUR; digit1<=ONE; digit2<=TWO; digit3<=SEVEN; end
      16'd7215: begin digit0<=FIVE; digit1<=ONE; digit2<=TWO; digit3<=SEVEN; end
      16'd7216: begin digit0<=SIX; digit1<=ONE; digit2<=TWO; digit3<=SEVEN; end
      16'd7217: begin digit0<=SEVEN; digit1<=ONE; digit2<=TWO; digit3<=SEVEN; end
      16'd7218: begin digit0<=EIGHT; digit1<=ONE; digit2<=TWO; digit3<=SEVEN; end
      16'd7219: begin digit0<=NINE; digit1<=ONE; digit2<=TWO; digit3<=SEVEN; end
      16'd7220: begin digit0<=ZERO; digit1<=TWO; digit2<=TWO; digit3<=SEVEN; end
      16'd7221: begin digit0<=ONE; digit1<=TWO; digit2<=TWO; digit3<=SEVEN; end
      16'd7222: begin digit0<=TWO; digit1<=TWO; digit2<=TWO; digit3<=SEVEN; end
      16'd7223: begin digit0<=THREE; digit1<=TWO; digit2<=TWO; digit3<=SEVEN; end
      16'd7224: begin digit0<=FOUR; digit1<=TWO; digit2<=TWO; digit3<=SEVEN; end
      16'd7225: begin digit0<=FIVE; digit1<=TWO; digit2<=TWO; digit3<=SEVEN; end
      16'd7226: begin digit0<=SIX; digit1<=TWO; digit2<=TWO; digit3<=SEVEN; end
      16'd7227: begin digit0<=SEVEN; digit1<=TWO; digit2<=TWO; digit3<=SEVEN; end
      16'd7228: begin digit0<=EIGHT; digit1<=TWO; digit2<=TWO; digit3<=SEVEN; end
      16'd7229: begin digit0<=NINE; digit1<=TWO; digit2<=TWO; digit3<=SEVEN; end
      16'd7230: begin digit0<=ZERO; digit1<=THREE; digit2<=TWO; digit3<=SEVEN; end
      16'd7231: begin digit0<=ONE; digit1<=THREE; digit2<=TWO; digit3<=SEVEN; end
      16'd7232: begin digit0<=TWO; digit1<=THREE; digit2<=TWO; digit3<=SEVEN; end
      16'd7233: begin digit0<=THREE; digit1<=THREE; digit2<=TWO; digit3<=SEVEN; end
      16'd7234: begin digit0<=FOUR; digit1<=THREE; digit2<=TWO; digit3<=SEVEN; end
      16'd7235: begin digit0<=FIVE; digit1<=THREE; digit2<=TWO; digit3<=SEVEN; end
      16'd7236: begin digit0<=SIX; digit1<=THREE; digit2<=TWO; digit3<=SEVEN; end
      16'd7237: begin digit0<=SEVEN; digit1<=THREE; digit2<=TWO; digit3<=SEVEN; end
      16'd7238: begin digit0<=EIGHT; digit1<=THREE; digit2<=TWO; digit3<=SEVEN; end
      16'd7239: begin digit0<=NINE; digit1<=THREE; digit2<=TWO; digit3<=SEVEN; end
      16'd7240: begin digit0<=ZERO; digit1<=FOUR; digit2<=TWO; digit3<=SEVEN; end
      16'd7241: begin digit0<=ONE; digit1<=FOUR; digit2<=TWO; digit3<=SEVEN; end
      16'd7242: begin digit0<=TWO; digit1<=FOUR; digit2<=TWO; digit3<=SEVEN; end
      16'd7243: begin digit0<=THREE; digit1<=FOUR; digit2<=TWO; digit3<=SEVEN; end
      16'd7244: begin digit0<=FOUR; digit1<=FOUR; digit2<=TWO; digit3<=SEVEN; end
      16'd7245: begin digit0<=FIVE; digit1<=FOUR; digit2<=TWO; digit3<=SEVEN; end
      16'd7246: begin digit0<=SIX; digit1<=FOUR; digit2<=TWO; digit3<=SEVEN; end
      16'd7247: begin digit0<=SEVEN; digit1<=FOUR; digit2<=TWO; digit3<=SEVEN; end
      16'd7248: begin digit0<=EIGHT; digit1<=FOUR; digit2<=TWO; digit3<=SEVEN; end
      16'd7249: begin digit0<=NINE; digit1<=FOUR; digit2<=TWO; digit3<=SEVEN; end
      16'd7250: begin digit0<=ZERO; digit1<=FIVE; digit2<=TWO; digit3<=SEVEN; end
      16'd7251: begin digit0<=ONE; digit1<=FIVE; digit2<=TWO; digit3<=SEVEN; end
      16'd7252: begin digit0<=TWO; digit1<=FIVE; digit2<=TWO; digit3<=SEVEN; end
      16'd7253: begin digit0<=THREE; digit1<=FIVE; digit2<=TWO; digit3<=SEVEN; end
      16'd7254: begin digit0<=FOUR; digit1<=FIVE; digit2<=TWO; digit3<=SEVEN; end
      16'd7255: begin digit0<=FIVE; digit1<=FIVE; digit2<=TWO; digit3<=SEVEN; end
      16'd7256: begin digit0<=SIX; digit1<=FIVE; digit2<=TWO; digit3<=SEVEN; end
      16'd7257: begin digit0<=SEVEN; digit1<=FIVE; digit2<=TWO; digit3<=SEVEN; end
      16'd7258: begin digit0<=EIGHT; digit1<=FIVE; digit2<=TWO; digit3<=SEVEN; end
      16'd7259: begin digit0<=NINE; digit1<=FIVE; digit2<=TWO; digit3<=SEVEN; end
      16'd7260: begin digit0<=ZERO; digit1<=SIX; digit2<=TWO; digit3<=SEVEN; end
      16'd7261: begin digit0<=ONE; digit1<=SIX; digit2<=TWO; digit3<=SEVEN; end
      16'd7262: begin digit0<=TWO; digit1<=SIX; digit2<=TWO; digit3<=SEVEN; end
      16'd7263: begin digit0<=THREE; digit1<=SIX; digit2<=TWO; digit3<=SEVEN; end
      16'd7264: begin digit0<=FOUR; digit1<=SIX; digit2<=TWO; digit3<=SEVEN; end
      16'd7265: begin digit0<=FIVE; digit1<=SIX; digit2<=TWO; digit3<=SEVEN; end
      16'd7266: begin digit0<=SIX; digit1<=SIX; digit2<=TWO; digit3<=SEVEN; end
      16'd7267: begin digit0<=SEVEN; digit1<=SIX; digit2<=TWO; digit3<=SEVEN; end
      16'd7268: begin digit0<=EIGHT; digit1<=SIX; digit2<=TWO; digit3<=SEVEN; end
      16'd7269: begin digit0<=NINE; digit1<=SIX; digit2<=TWO; digit3<=SEVEN; end
      16'd7270: begin digit0<=ZERO; digit1<=SEVEN; digit2<=TWO; digit3<=SEVEN; end
      16'd7271: begin digit0<=ONE; digit1<=SEVEN; digit2<=TWO; digit3<=SEVEN; end
      16'd7272: begin digit0<=TWO; digit1<=SEVEN; digit2<=TWO; digit3<=SEVEN; end
      16'd7273: begin digit0<=THREE; digit1<=SEVEN; digit2<=TWO; digit3<=SEVEN; end
      16'd7274: begin digit0<=FOUR; digit1<=SEVEN; digit2<=TWO; digit3<=SEVEN; end
      16'd7275: begin digit0<=FIVE; digit1<=SEVEN; digit2<=TWO; digit3<=SEVEN; end
      16'd7276: begin digit0<=SIX; digit1<=SEVEN; digit2<=TWO; digit3<=SEVEN; end
      16'd7277: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=TWO; digit3<=SEVEN; end
      16'd7278: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=TWO; digit3<=SEVEN; end
      16'd7279: begin digit0<=NINE; digit1<=SEVEN; digit2<=TWO; digit3<=SEVEN; end
      16'd7280: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=SEVEN; end
      16'd7281: begin digit0<=ONE; digit1<=EIGHT; digit2<=TWO; digit3<=SEVEN; end
      16'd7282: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=SEVEN; end
      16'd7283: begin digit0<=THREE; digit1<=EIGHT; digit2<=TWO; digit3<=SEVEN; end
      16'd7284: begin digit0<=FOUR; digit1<=EIGHT; digit2<=TWO; digit3<=SEVEN; end
      16'd7285: begin digit0<=FIVE; digit1<=EIGHT; digit2<=TWO; digit3<=SEVEN; end
      16'd7286: begin digit0<=SIX; digit1<=EIGHT; digit2<=TWO; digit3<=SEVEN; end
      16'd7287: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=TWO; digit3<=SEVEN; end
      16'd7288: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=TWO; digit3<=SEVEN; end
      16'd7289: begin digit0<=NINE; digit1<=EIGHT; digit2<=TWO; digit3<=SEVEN; end
      16'd7290: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=SEVEN; end
      16'd7291: begin digit0<=ONE; digit1<=NINE; digit2<=TWO; digit3<=SEVEN; end
      16'd7292: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=SEVEN; end
      16'd7293: begin digit0<=THREE; digit1<=NINE; digit2<=TWO; digit3<=SEVEN; end
      16'd7294: begin digit0<=FOUR; digit1<=NINE; digit2<=TWO; digit3<=SEVEN; end
      16'd7295: begin digit0<=FIVE; digit1<=NINE; digit2<=TWO; digit3<=SEVEN; end
      16'd7296: begin digit0<=SIX; digit1<=NINE; digit2<=TWO; digit3<=SEVEN; end
      16'd7297: begin digit0<=SEVEN; digit1<=NINE; digit2<=TWO; digit3<=SEVEN; end
      16'd7298: begin digit0<=EIGHT; digit1<=NINE; digit2<=TWO; digit3<=SEVEN; end
      16'd7299: begin digit0<=NINE; digit1<=NINE; digit2<=TWO; digit3<=SEVEN; end
	  16'd7300: begin digit0<=ZERO; digit1<=ZERO; digit2<=THREE; digit3<=SEVEN; end
      16'd7301: begin digit0<=ONE; digit1<=ZERO; digit2<=THREE; digit3<=SEVEN; end
      16'd7302: begin digit0<=TWO; digit1<=ZERO; digit2<=THREE; digit3<=SEVEN; end
      16'd7303: begin digit0<=THREE; digit1<=ZERO; digit2<=THREE; digit3<=SEVEN; end
      16'd7304: begin digit0<=FOUR; digit1<=ZERO; digit2<=THREE; digit3<=SEVEN; end
      16'd7305: begin digit0<=FIVE; digit1<=ZERO; digit2<=THREE; digit3<=SEVEN; end
      16'd7306: begin digit0<=SIX; digit1<=ZERO; digit2<=THREE; digit3<=SEVEN; end
      16'd7307: begin digit0<=SEVEN; digit1<=ZERO; digit2<=THREE; digit3<=SEVEN; end
      16'd7308: begin digit0<=EIGHT; digit1<=ZERO; digit2<=THREE; digit3<=SEVEN; end
      16'd7309: begin digit0<=NINE; digit1<=ZERO; digit2<=THREE; digit3<=SEVEN; end
      16'd7310: begin digit0<=ZERO; digit1<=ONE; digit2<=THREE; digit3<=SEVEN; end
      16'd7311: begin digit0<=ONE; digit1<=ONE; digit2<=THREE; digit3<=SEVEN; end
      16'd7312: begin digit0<=TWO; digit1<=ONE; digit2<=THREE; digit3<=SEVEN; end
      16'd7313: begin digit0<=THREE; digit1<=ONE; digit2<=THREE; digit3<=SEVEN; end
      16'd7314: begin digit0<=FOUR; digit1<=ONE; digit2<=THREE; digit3<=SEVEN; end
      16'd7315: begin digit0<=FIVE; digit1<=ONE; digit2<=THREE; digit3<=SEVEN; end
      16'd7316: begin digit0<=SIX; digit1<=ONE; digit2<=THREE; digit3<=SEVEN; end
      16'd7317: begin digit0<=SEVEN; digit1<=ONE; digit2<=THREE; digit3<=SEVEN; end
      16'd7318: begin digit0<=EIGHT; digit1<=ONE; digit2<=THREE; digit3<=SEVEN; end
      16'd7319: begin digit0<=NINE; digit1<=ONE; digit2<=THREE; digit3<=SEVEN; end
      16'd7320: begin digit0<=ZERO; digit1<=TWO; digit2<=THREE; digit3<=SEVEN; end
      16'd7321: begin digit0<=ONE; digit1<=TWO; digit2<=THREE; digit3<=SEVEN; end
      16'd7322: begin digit0<=TWO; digit1<=TWO; digit2<=THREE; digit3<=SEVEN; end
      16'd7323: begin digit0<=THREE; digit1<=TWO; digit2<=THREE; digit3<=SEVEN; end
      16'd7324: begin digit0<=FOUR; digit1<=TWO; digit2<=THREE; digit3<=SEVEN; end
      16'd7325: begin digit0<=FIVE; digit1<=TWO; digit2<=THREE; digit3<=SEVEN; end
      16'd7326: begin digit0<=SIX; digit1<=TWO; digit2<=THREE; digit3<=SEVEN; end
      16'd7327: begin digit0<=SEVEN; digit1<=TWO; digit2<=THREE; digit3<=SEVEN; end
      16'd7328: begin digit0<=EIGHT; digit1<=TWO; digit2<=THREE; digit3<=SEVEN; end
      16'd7329: begin digit0<=NINE; digit1<=TWO; digit2<=THREE; digit3<=SEVEN; end
      16'd7330: begin digit0<=ZERO; digit1<=THREE; digit2<=THREE; digit3<=SEVEN; end
      16'd7331: begin digit0<=ONE; digit1<=THREE; digit2<=THREE; digit3<=SEVEN; end
      16'd7332: begin digit0<=TWO; digit1<=THREE; digit2<=THREE; digit3<=SEVEN; end
      16'd7333: begin digit0<=THREE; digit1<=THREE; digit2<=THREE; digit3<=SEVEN; end
      16'd7334: begin digit0<=FOUR; digit1<=THREE; digit2<=THREE; digit3<=SEVEN; end
      16'd7335: begin digit0<=FIVE; digit1<=THREE; digit2<=THREE; digit3<=SEVEN; end
      16'd7336: begin digit0<=SIX; digit1<=THREE; digit2<=THREE; digit3<=SEVEN; end
      16'd7337: begin digit0<=SEVEN; digit1<=THREE; digit2<=THREE; digit3<=SEVEN; end
      16'd7338: begin digit0<=EIGHT; digit1<=THREE; digit2<=THREE; digit3<=SEVEN; end
      16'd7339: begin digit0<=NINE; digit1<=THREE; digit2<=THREE; digit3<=SEVEN; end
      16'd7340: begin digit0<=ZERO; digit1<=FOUR; digit2<=THREE; digit3<=SEVEN; end
      16'd7341: begin digit0<=ONE; digit1<=FOUR; digit2<=THREE; digit3<=SEVEN; end
      16'd7342: begin digit0<=TWO; digit1<=FOUR; digit2<=THREE; digit3<=SEVEN; end
      16'd7343: begin digit0<=THREE; digit1<=FOUR; digit2<=THREE; digit3<=SEVEN; end
      16'd7344: begin digit0<=FOUR; digit1<=FOUR; digit2<=THREE; digit3<=SEVEN; end
      16'd7345: begin digit0<=FIVE; digit1<=FOUR; digit2<=THREE; digit3<=SEVEN; end
      16'd7346: begin digit0<=SIX; digit1<=FOUR; digit2<=THREE; digit3<=SEVEN; end
      16'd7347: begin digit0<=SEVEN; digit1<=FOUR; digit2<=THREE; digit3<=SEVEN; end
      16'd7348: begin digit0<=EIGHT; digit1<=FOUR; digit2<=THREE; digit3<=SEVEN; end
      16'd7349: begin digit0<=NINE; digit1<=FOUR; digit2<=THREE; digit3<=SEVEN; end
      16'd7350: begin digit0<=ZERO; digit1<=FIVE; digit2<=THREE; digit3<=SEVEN; end
      16'd7351: begin digit0<=ONE; digit1<=FIVE; digit2<=THREE; digit3<=SEVEN; end
      16'd7352: begin digit0<=TWO; digit1<=FIVE; digit2<=THREE; digit3<=SEVEN; end
      16'd7353: begin digit0<=THREE; digit1<=FIVE; digit2<=THREE; digit3<=SEVEN; end
      16'd7354: begin digit0<=FOUR; digit1<=FIVE; digit2<=THREE; digit3<=SEVEN; end
      16'd7355: begin digit0<=FIVE; digit1<=FIVE; digit2<=THREE; digit3<=SEVEN; end
      16'd7356: begin digit0<=SIX; digit1<=FIVE; digit2<=THREE; digit3<=SEVEN; end
      16'd7357: begin digit0<=SEVEN; digit1<=FIVE; digit2<=THREE; digit3<=SEVEN; end
      16'd7358: begin digit0<=EIGHT; digit1<=FIVE; digit2<=THREE; digit3<=SEVEN; end
      16'd7359: begin digit0<=NINE; digit1<=FIVE; digit2<=THREE; digit3<=SEVEN; end
      16'd7360: begin digit0<=ZERO; digit1<=SIX; digit2<=THREE; digit3<=SEVEN; end
      16'd7361: begin digit0<=ONE; digit1<=SIX; digit2<=THREE; digit3<=SEVEN; end
      16'd7362: begin digit0<=TWO; digit1<=SIX; digit2<=THREE; digit3<=SEVEN; end
      16'd7363: begin digit0<=THREE; digit1<=SIX; digit2<=THREE; digit3<=SEVEN; end
      16'd7364: begin digit0<=FOUR; digit1<=SIX; digit2<=THREE; digit3<=SEVEN; end
      16'd7365: begin digit0<=FIVE; digit1<=SIX; digit2<=THREE; digit3<=SEVEN; end
      16'd7366: begin digit0<=SIX; digit1<=SIX; digit2<=THREE; digit3<=SEVEN; end
      16'd7367: begin digit0<=SEVEN; digit1<=SIX; digit2<=THREE; digit3<=SEVEN; end
      16'd7368: begin digit0<=EIGHT; digit1<=SIX; digit2<=THREE; digit3<=SEVEN; end
      16'd7369: begin digit0<=NINE; digit1<=SIX; digit2<=THREE; digit3<=SEVEN; end
      16'd7370: begin digit0<=ZERO; digit1<=SEVEN; digit2<=THREE; digit3<=SEVEN; end
      16'd7371: begin digit0<=ONE; digit1<=SEVEN; digit2<=THREE; digit3<=SEVEN; end
      16'd7372: begin digit0<=TWO; digit1<=SEVEN; digit2<=THREE; digit3<=SEVEN; end
      16'd7373: begin digit0<=THREE; digit1<=SEVEN; digit2<=THREE; digit3<=SEVEN; end
      16'd7374: begin digit0<=FOUR; digit1<=SEVEN; digit2<=THREE; digit3<=SEVEN; end
      16'd7375: begin digit0<=FIVE; digit1<=SEVEN; digit2<=THREE; digit3<=SEVEN; end
      16'd7376: begin digit0<=SIX; digit1<=SEVEN; digit2<=THREE; digit3<=SEVEN; end
      16'd7377: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=THREE; digit3<=SEVEN; end
      16'd7378: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=THREE; digit3<=SEVEN; end
      16'd7379: begin digit0<=NINE; digit1<=SEVEN; digit2<=THREE; digit3<=SEVEN; end
      16'd7380: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=SEVEN; end
      16'd7381: begin digit0<=ONE; digit1<=EIGHT; digit2<=THREE; digit3<=SEVEN; end
      16'd7382: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=SEVEN; end
      16'd7383: begin digit0<=THREE; digit1<=EIGHT; digit2<=THREE; digit3<=SEVEN; end
      16'd7384: begin digit0<=FOUR; digit1<=EIGHT; digit2<=THREE; digit3<=SEVEN; end
      16'd7385: begin digit0<=FIVE; digit1<=EIGHT; digit2<=THREE; digit3<=SEVEN; end
      16'd7386: begin digit0<=SIX; digit1<=EIGHT; digit2<=THREE; digit3<=SEVEN; end
      16'd7387: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=THREE; digit3<=SEVEN; end
      16'd7388: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=THREE; digit3<=SEVEN; end
      16'd7389: begin digit0<=NINE; digit1<=EIGHT; digit2<=THREE; digit3<=SEVEN; end
      16'd7390: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=SEVEN; end
      16'd7391: begin digit0<=ONE; digit1<=NINE; digit2<=THREE; digit3<=SEVEN; end
      16'd7392: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=SEVEN; end
      16'd7393: begin digit0<=THREE; digit1<=NINE; digit2<=THREE; digit3<=SEVEN; end
      16'd7394: begin digit0<=FOUR; digit1<=NINE; digit2<=THREE; digit3<=SEVEN; end
      16'd7395: begin digit0<=FIVE; digit1<=NINE; digit2<=THREE; digit3<=SEVEN; end
      16'd7396: begin digit0<=SIX; digit1<=NINE; digit2<=THREE; digit3<=SEVEN; end
      16'd7397: begin digit0<=SEVEN; digit1<=NINE; digit2<=THREE; digit3<=SEVEN; end
      16'd7398: begin digit0<=EIGHT; digit1<=NINE; digit2<=THREE; digit3<=SEVEN; end
      16'd7399: begin digit0<=NINE; digit1<=NINE; digit2<=THREE; digit3<=SEVEN; end
	  16'd7400: begin digit0<=ZERO; digit1<=ZERO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7401: begin digit0<=ONE; digit1<=ZERO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7402: begin digit0<=TWO; digit1<=ZERO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7403: begin digit0<=THREE; digit1<=ZERO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7404: begin digit0<=FOUR; digit1<=ZERO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7405: begin digit0<=FIVE; digit1<=ZERO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7406: begin digit0<=SIX; digit1<=ZERO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7407: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7408: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7409: begin digit0<=NINE; digit1<=ZERO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7410: begin digit0<=ZERO; digit1<=ONE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7411: begin digit0<=ONE; digit1<=ONE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7412: begin digit0<=TWO; digit1<=ONE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7413: begin digit0<=THREE; digit1<=ONE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7414: begin digit0<=FOUR; digit1<=ONE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7415: begin digit0<=FIVE; digit1<=ONE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7416: begin digit0<=SIX; digit1<=ONE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7417: begin digit0<=SEVEN; digit1<=ONE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7418: begin digit0<=EIGHT; digit1<=ONE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7419: begin digit0<=NINE; digit1<=ONE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7420: begin digit0<=ZERO; digit1<=TWO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7421: begin digit0<=ONE; digit1<=TWO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7422: begin digit0<=TWO; digit1<=TWO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7423: begin digit0<=THREE; digit1<=TWO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7424: begin digit0<=FOUR; digit1<=TWO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7425: begin digit0<=FIVE; digit1<=TWO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7426: begin digit0<=SIX; digit1<=TWO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7427: begin digit0<=SEVEN; digit1<=TWO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7428: begin digit0<=EIGHT; digit1<=TWO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7429: begin digit0<=NINE; digit1<=TWO; digit2<=FOUR; digit3<=SEVEN; end
      16'd7430: begin digit0<=ZERO; digit1<=THREE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7431: begin digit0<=ONE; digit1<=THREE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7432: begin digit0<=TWO; digit1<=THREE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7433: begin digit0<=THREE; digit1<=THREE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7434: begin digit0<=FOUR; digit1<=THREE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7435: begin digit0<=FIVE; digit1<=THREE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7436: begin digit0<=SIX; digit1<=THREE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7437: begin digit0<=SEVEN; digit1<=THREE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7438: begin digit0<=EIGHT; digit1<=THREE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7439: begin digit0<=NINE; digit1<=THREE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7440: begin digit0<=ZERO; digit1<=FOUR; digit2<=FOUR; digit3<=SEVEN; end
      16'd7441: begin digit0<=ONE; digit1<=FOUR; digit2<=FOUR; digit3<=SEVEN; end
      16'd7442: begin digit0<=TWO; digit1<=FOUR; digit2<=FOUR; digit3<=SEVEN; end
      16'd7443: begin digit0<=THREE; digit1<=FOUR; digit2<=FOUR; digit3<=SEVEN; end
      16'd7444: begin digit0<=FOUR; digit1<=FOUR; digit2<=FOUR; digit3<=SEVEN; end
      16'd7445: begin digit0<=FIVE; digit1<=FOUR; digit2<=FOUR; digit3<=SEVEN; end
      16'd7446: begin digit0<=SIX; digit1<=FOUR; digit2<=FOUR; digit3<=SEVEN; end
      16'd7447: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FOUR; digit3<=SEVEN; end
      16'd7448: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FOUR; digit3<=SEVEN; end
      16'd7449: begin digit0<=NINE; digit1<=FOUR; digit2<=FOUR; digit3<=SEVEN; end
      16'd7450: begin digit0<=ZERO; digit1<=FIVE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7451: begin digit0<=ONE; digit1<=FIVE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7452: begin digit0<=TWO; digit1<=FIVE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7453: begin digit0<=THREE; digit1<=FIVE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7454: begin digit0<=FOUR; digit1<=FIVE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7455: begin digit0<=FIVE; digit1<=FIVE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7456: begin digit0<=SIX; digit1<=FIVE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7457: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7458: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7459: begin digit0<=NINE; digit1<=FIVE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7460: begin digit0<=ZERO; digit1<=SIX; digit2<=FOUR; digit3<=SEVEN; end
      16'd7461: begin digit0<=ONE; digit1<=SIX; digit2<=FOUR; digit3<=SEVEN; end
      16'd7462: begin digit0<=TWO; digit1<=SIX; digit2<=FOUR; digit3<=SEVEN; end
      16'd7463: begin digit0<=THREE; digit1<=SIX; digit2<=FOUR; digit3<=SEVEN; end
      16'd7464: begin digit0<=FOUR; digit1<=SIX; digit2<=FOUR; digit3<=SEVEN; end
      16'd7465: begin digit0<=FIVE; digit1<=SIX; digit2<=FOUR; digit3<=SEVEN; end
      16'd7466: begin digit0<=SIX; digit1<=SIX; digit2<=FOUR; digit3<=SEVEN; end
      16'd7467: begin digit0<=SEVEN; digit1<=SIX; digit2<=FOUR; digit3<=SEVEN; end
      16'd7468: begin digit0<=EIGHT; digit1<=SIX; digit2<=FOUR; digit3<=SEVEN; end
      16'd7469: begin digit0<=NINE; digit1<=SIX; digit2<=FOUR; digit3<=SEVEN; end
      16'd7470: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FOUR; digit3<=SEVEN; end
      16'd7471: begin digit0<=ONE; digit1<=SEVEN; digit2<=FOUR; digit3<=SEVEN; end
      16'd7472: begin digit0<=TWO; digit1<=SEVEN; digit2<=FOUR; digit3<=SEVEN; end
      16'd7473: begin digit0<=THREE; digit1<=SEVEN; digit2<=FOUR; digit3<=SEVEN; end
      16'd7474: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FOUR; digit3<=SEVEN; end
      16'd7475: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FOUR; digit3<=SEVEN; end
      16'd7476: begin digit0<=SIX; digit1<=SEVEN; digit2<=FOUR; digit3<=SEVEN; end
      16'd7477: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FOUR; digit3<=SEVEN; end
      16'd7478: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FOUR; digit3<=SEVEN; end
      16'd7479: begin digit0<=NINE; digit1<=SEVEN; digit2<=FOUR; digit3<=SEVEN; end
      16'd7480: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=SEVEN; end
      16'd7481: begin digit0<=ONE; digit1<=EIGHT; digit2<=FOUR; digit3<=SEVEN; end
      16'd7482: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=SEVEN; end
      16'd7483: begin digit0<=THREE; digit1<=EIGHT; digit2<=FOUR; digit3<=SEVEN; end
      16'd7484: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FOUR; digit3<=SEVEN; end
      16'd7485: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FOUR; digit3<=SEVEN; end
      16'd7486: begin digit0<=SIX; digit1<=EIGHT; digit2<=FOUR; digit3<=SEVEN; end
      16'd7487: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FOUR; digit3<=SEVEN; end
      16'd7488: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FOUR; digit3<=SEVEN; end
      16'd7489: begin digit0<=NINE; digit1<=EIGHT; digit2<=FOUR; digit3<=SEVEN; end
      16'd7490: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7491: begin digit0<=ONE; digit1<=NINE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7492: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7493: begin digit0<=THREE; digit1<=NINE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7494: begin digit0<=FOUR; digit1<=NINE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7495: begin digit0<=FIVE; digit1<=NINE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7496: begin digit0<=SIX; digit1<=NINE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7497: begin digit0<=SEVEN; digit1<=NINE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7498: begin digit0<=EIGHT; digit1<=NINE; digit2<=FOUR; digit3<=SEVEN; end
      16'd7499: begin digit0<=NINE; digit1<=NINE; digit2<=FOUR; digit3<=SEVEN; end
	  16'd7500: begin digit0<=ZERO; digit1<=ZERO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7501: begin digit0<=ONE; digit1<=ZERO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7502: begin digit0<=TWO; digit1<=ZERO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7503: begin digit0<=THREE; digit1<=ZERO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7504: begin digit0<=FOUR; digit1<=ZERO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7505: begin digit0<=FIVE; digit1<=ZERO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7506: begin digit0<=SIX; digit1<=ZERO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7507: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7508: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7509: begin digit0<=NINE; digit1<=ZERO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7510: begin digit0<=ZERO; digit1<=ONE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7511: begin digit0<=ONE; digit1<=ONE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7512: begin digit0<=TWO; digit1<=ONE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7513: begin digit0<=THREE; digit1<=ONE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7514: begin digit0<=FOUR; digit1<=ONE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7515: begin digit0<=FIVE; digit1<=ONE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7516: begin digit0<=SIX; digit1<=ONE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7517: begin digit0<=SEVEN; digit1<=ONE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7518: begin digit0<=EIGHT; digit1<=ONE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7519: begin digit0<=NINE; digit1<=ONE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7520: begin digit0<=ZERO; digit1<=TWO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7521: begin digit0<=ONE; digit1<=TWO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7522: begin digit0<=TWO; digit1<=TWO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7523: begin digit0<=THREE; digit1<=TWO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7524: begin digit0<=FOUR; digit1<=TWO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7525: begin digit0<=FIVE; digit1<=TWO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7526: begin digit0<=SIX; digit1<=TWO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7527: begin digit0<=SEVEN; digit1<=TWO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7528: begin digit0<=EIGHT; digit1<=TWO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7529: begin digit0<=NINE; digit1<=TWO; digit2<=FIVE; digit3<=SEVEN; end
      16'd7530: begin digit0<=ZERO; digit1<=THREE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7531: begin digit0<=ONE; digit1<=THREE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7532: begin digit0<=TWO; digit1<=THREE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7533: begin digit0<=THREE; digit1<=THREE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7534: begin digit0<=FOUR; digit1<=THREE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7535: begin digit0<=FIVE; digit1<=THREE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7536: begin digit0<=SIX; digit1<=THREE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7537: begin digit0<=SEVEN; digit1<=THREE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7538: begin digit0<=EIGHT; digit1<=THREE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7539: begin digit0<=NINE; digit1<=THREE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7540: begin digit0<=ZERO; digit1<=FOUR; digit2<=FIVE; digit3<=SEVEN; end
      16'd7541: begin digit0<=ONE; digit1<=FOUR; digit2<=FIVE; digit3<=SEVEN; end
      16'd7542: begin digit0<=TWO; digit1<=FOUR; digit2<=FIVE; digit3<=SEVEN; end
      16'd7543: begin digit0<=THREE; digit1<=FOUR; digit2<=FIVE; digit3<=SEVEN; end
      16'd7544: begin digit0<=FOUR; digit1<=FOUR; digit2<=FIVE; digit3<=SEVEN; end
      16'd7545: begin digit0<=FIVE; digit1<=FOUR; digit2<=FIVE; digit3<=SEVEN; end
      16'd7546: begin digit0<=SIX; digit1<=FOUR; digit2<=FIVE; digit3<=SEVEN; end
      16'd7547: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FIVE; digit3<=SEVEN; end
      16'd7548: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FIVE; digit3<=SEVEN; end
      16'd7549: begin digit0<=NINE; digit1<=FOUR; digit2<=FIVE; digit3<=SEVEN; end
      16'd7550: begin digit0<=ZERO; digit1<=FIVE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7551: begin digit0<=ONE; digit1<=FIVE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7552: begin digit0<=TWO; digit1<=FIVE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7553: begin digit0<=THREE; digit1<=FIVE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7554: begin digit0<=FOUR; digit1<=FIVE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7555: begin digit0<=FIVE; digit1<=FIVE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7556: begin digit0<=SIX; digit1<=FIVE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7557: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7558: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7559: begin digit0<=NINE; digit1<=FIVE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7560: begin digit0<=ZERO; digit1<=SIX; digit2<=FIVE; digit3<=SEVEN; end
      16'd7561: begin digit0<=ONE; digit1<=SIX; digit2<=FIVE; digit3<=SEVEN; end
      16'd7562: begin digit0<=TWO; digit1<=SIX; digit2<=FIVE; digit3<=SEVEN; end
      16'd7563: begin digit0<=THREE; digit1<=SIX; digit2<=FIVE; digit3<=SEVEN; end
      16'd7564: begin digit0<=FOUR; digit1<=SIX; digit2<=FIVE; digit3<=SEVEN; end
      16'd7565: begin digit0<=FIVE; digit1<=SIX; digit2<=FIVE; digit3<=SEVEN; end
      16'd7566: begin digit0<=SIX; digit1<=SIX; digit2<=FIVE; digit3<=SEVEN; end
      16'd7567: begin digit0<=SEVEN; digit1<=SIX; digit2<=FIVE; digit3<=SEVEN; end
      16'd7568: begin digit0<=EIGHT; digit1<=SIX; digit2<=FIVE; digit3<=SEVEN; end
      16'd7569: begin digit0<=NINE; digit1<=SIX; digit2<=FIVE; digit3<=SEVEN; end
      16'd7570: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FIVE; digit3<=SEVEN; end
      16'd7571: begin digit0<=ONE; digit1<=SEVEN; digit2<=FIVE; digit3<=SEVEN; end
      16'd7572: begin digit0<=TWO; digit1<=SEVEN; digit2<=FIVE; digit3<=SEVEN; end
      16'd7573: begin digit0<=THREE; digit1<=SEVEN; digit2<=FIVE; digit3<=SEVEN; end
      16'd7574: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FIVE; digit3<=SEVEN; end
      16'd7575: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FIVE; digit3<=SEVEN; end
      16'd7576: begin digit0<=SIX; digit1<=SEVEN; digit2<=FIVE; digit3<=SEVEN; end
      16'd7577: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FIVE; digit3<=SEVEN; end
      16'd7578: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FIVE; digit3<=SEVEN; end
      16'd7579: begin digit0<=NINE; digit1<=SEVEN; digit2<=FIVE; digit3<=SEVEN; end
      16'd7580: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=SEVEN; end
      16'd7581: begin digit0<=ONE; digit1<=EIGHT; digit2<=FIVE; digit3<=SEVEN; end
      16'd7582: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=SEVEN; end
      16'd7583: begin digit0<=THREE; digit1<=EIGHT; digit2<=FIVE; digit3<=SEVEN; end
      16'd7584: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FIVE; digit3<=SEVEN; end
      16'd7585: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FIVE; digit3<=SEVEN; end
      16'd7586: begin digit0<=SIX; digit1<=EIGHT; digit2<=FIVE; digit3<=SEVEN; end
      16'd7587: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FIVE; digit3<=SEVEN; end
      16'd7588: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FIVE; digit3<=SEVEN; end
      16'd7589: begin digit0<=NINE; digit1<=EIGHT; digit2<=FIVE; digit3<=SEVEN; end
      16'd7590: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7591: begin digit0<=ONE; digit1<=NINE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7592: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7593: begin digit0<=THREE; digit1<=NINE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7594: begin digit0<=FOUR; digit1<=NINE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7595: begin digit0<=FIVE; digit1<=NINE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7596: begin digit0<=SIX; digit1<=NINE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7597: begin digit0<=SEVEN; digit1<=NINE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7598: begin digit0<=EIGHT; digit1<=NINE; digit2<=FIVE; digit3<=SEVEN; end
      16'd7599: begin digit0<=NINE; digit1<=NINE; digit2<=FIVE; digit3<=SEVEN; end
	  16'd7600: begin digit0<=ZERO; digit1<=ZERO; digit2<=SIX; digit3<=SEVEN; end
      16'd7601: begin digit0<=ONE; digit1<=ZERO; digit2<=SIX; digit3<=SEVEN; end
      16'd7602: begin digit0<=TWO; digit1<=ZERO; digit2<=SIX; digit3<=SEVEN; end
      16'd7603: begin digit0<=THREE; digit1<=ZERO; digit2<=SIX; digit3<=SEVEN; end
      16'd7604: begin digit0<=FOUR; digit1<=ZERO; digit2<=SIX; digit3<=SEVEN; end
      16'd7605: begin digit0<=FIVE; digit1<=ZERO; digit2<=SIX; digit3<=SEVEN; end
      16'd7606: begin digit0<=SIX; digit1<=ZERO; digit2<=SIX; digit3<=SEVEN; end
      16'd7607: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SIX; digit3<=SEVEN; end
      16'd7608: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SIX; digit3<=SEVEN; end
      16'd7609: begin digit0<=NINE; digit1<=ZERO; digit2<=SIX; digit3<=SEVEN; end
      16'd7610: begin digit0<=ZERO; digit1<=ONE; digit2<=SIX; digit3<=SEVEN; end
      16'd7611: begin digit0<=ONE; digit1<=ONE; digit2<=SIX; digit3<=SEVEN; end
      16'd7612: begin digit0<=TWO; digit1<=ONE; digit2<=SIX; digit3<=SEVEN; end
      16'd7613: begin digit0<=THREE; digit1<=ONE; digit2<=SIX; digit3<=SEVEN; end
      16'd7614: begin digit0<=FOUR; digit1<=ONE; digit2<=SIX; digit3<=SEVEN; end
      16'd7615: begin digit0<=FIVE; digit1<=ONE; digit2<=SIX; digit3<=SEVEN; end
      16'd7616: begin digit0<=SIX; digit1<=ONE; digit2<=SIX; digit3<=SEVEN; end
      16'd7617: begin digit0<=SEVEN; digit1<=ONE; digit2<=SIX; digit3<=SEVEN; end
      16'd7618: begin digit0<=EIGHT; digit1<=ONE; digit2<=SIX; digit3<=SEVEN; end
      16'd7619: begin digit0<=NINE; digit1<=ONE; digit2<=SIX; digit3<=SEVEN; end
      16'd7620: begin digit0<=ZERO; digit1<=TWO; digit2<=SIX; digit3<=SEVEN; end
      16'd7621: begin digit0<=ONE; digit1<=TWO; digit2<=SIX; digit3<=SEVEN; end
      16'd7622: begin digit0<=TWO; digit1<=TWO; digit2<=SIX; digit3<=SEVEN; end
      16'd7623: begin digit0<=THREE; digit1<=TWO; digit2<=SIX; digit3<=SEVEN; end
      16'd7624: begin digit0<=FOUR; digit1<=TWO; digit2<=SIX; digit3<=SEVEN; end
      16'd7625: begin digit0<=FIVE; digit1<=TWO; digit2<=SIX; digit3<=SEVEN; end
      16'd7626: begin digit0<=SIX; digit1<=TWO; digit2<=SIX; digit3<=SEVEN; end
      16'd7627: begin digit0<=SEVEN; digit1<=TWO; digit2<=SIX; digit3<=SEVEN; end
      16'd7628: begin digit0<=EIGHT; digit1<=TWO; digit2<=SIX; digit3<=SEVEN; end
      16'd7629: begin digit0<=NINE; digit1<=TWO; digit2<=SIX; digit3<=SEVEN; end
      16'd7630: begin digit0<=ZERO; digit1<=THREE; digit2<=SIX; digit3<=SEVEN; end
      16'd7631: begin digit0<=ONE; digit1<=THREE; digit2<=SIX; digit3<=SEVEN; end
      16'd7632: begin digit0<=TWO; digit1<=THREE; digit2<=SIX; digit3<=SEVEN; end
      16'd7633: begin digit0<=THREE; digit1<=THREE; digit2<=SIX; digit3<=SEVEN; end
      16'd7634: begin digit0<=FOUR; digit1<=THREE; digit2<=SIX; digit3<=SEVEN; end
      16'd7635: begin digit0<=FIVE; digit1<=THREE; digit2<=SIX; digit3<=SEVEN; end
      16'd7636: begin digit0<=SIX; digit1<=THREE; digit2<=SIX; digit3<=SEVEN; end
      16'd7637: begin digit0<=SEVEN; digit1<=THREE; digit2<=SIX; digit3<=SEVEN; end
      16'd7638: begin digit0<=EIGHT; digit1<=THREE; digit2<=SIX; digit3<=SEVEN; end
      16'd7639: begin digit0<=NINE; digit1<=THREE; digit2<=SIX; digit3<=SEVEN; end
      16'd7640: begin digit0<=ZERO; digit1<=FOUR; digit2<=SIX; digit3<=SEVEN; end
      16'd7641: begin digit0<=ONE; digit1<=FOUR; digit2<=SIX; digit3<=SEVEN; end
      16'd7642: begin digit0<=TWO; digit1<=FOUR; digit2<=SIX; digit3<=SEVEN; end
      16'd7643: begin digit0<=THREE; digit1<=FOUR; digit2<=SIX; digit3<=SEVEN; end
      16'd7644: begin digit0<=FOUR; digit1<=FOUR; digit2<=SIX; digit3<=SEVEN; end
      16'd7645: begin digit0<=FIVE; digit1<=FOUR; digit2<=SIX; digit3<=SEVEN; end
      16'd7646: begin digit0<=SIX; digit1<=FOUR; digit2<=SIX; digit3<=SEVEN; end
      16'd7647: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SIX; digit3<=SEVEN; end
      16'd7648: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SIX; digit3<=SEVEN; end
      16'd7649: begin digit0<=NINE; digit1<=FOUR; digit2<=SIX; digit3<=SEVEN; end
      16'd7650: begin digit0<=ZERO; digit1<=FIVE; digit2<=SIX; digit3<=SEVEN; end
      16'd7651: begin digit0<=ONE; digit1<=FIVE; digit2<=SIX; digit3<=SEVEN; end
      16'd7652: begin digit0<=TWO; digit1<=FIVE; digit2<=SIX; digit3<=SEVEN; end
      16'd7653: begin digit0<=THREE; digit1<=FIVE; digit2<=SIX; digit3<=SEVEN; end
      16'd7654: begin digit0<=FOUR; digit1<=FIVE; digit2<=SIX; digit3<=SEVEN; end
      16'd7655: begin digit0<=FIVE; digit1<=FIVE; digit2<=SIX; digit3<=SEVEN; end
      16'd7656: begin digit0<=SIX; digit1<=FIVE; digit2<=SIX; digit3<=SEVEN; end
      16'd7657: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SIX; digit3<=SEVEN; end
      16'd7658: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SIX; digit3<=SEVEN; end
      16'd7659: begin digit0<=NINE; digit1<=FIVE; digit2<=SIX; digit3<=SEVEN; end
      16'd7660: begin digit0<=ZERO; digit1<=SIX; digit2<=SIX; digit3<=SEVEN; end
      16'd7661: begin digit0<=ONE; digit1<=SIX; digit2<=SIX; digit3<=SEVEN; end
      16'd7662: begin digit0<=TWO; digit1<=SIX; digit2<=SIX; digit3<=SEVEN; end
      16'd7663: begin digit0<=THREE; digit1<=SIX; digit2<=SIX; digit3<=SEVEN; end
      16'd7664: begin digit0<=FOUR; digit1<=SIX; digit2<=SIX; digit3<=SEVEN; end
      16'd7665: begin digit0<=FIVE; digit1<=SIX; digit2<=SIX; digit3<=SEVEN; end
      16'd7666: begin digit0<=SIX; digit1<=SIX; digit2<=SIX; digit3<=SEVEN; end
      16'd7667: begin digit0<=SEVEN; digit1<=SIX; digit2<=SIX; digit3<=SEVEN; end
      16'd7668: begin digit0<=EIGHT; digit1<=SIX; digit2<=SIX; digit3<=SEVEN; end
      16'd7669: begin digit0<=NINE; digit1<=SIX; digit2<=SIX; digit3<=SEVEN; end
      16'd7670: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SIX; digit3<=SEVEN; end
      16'd7671: begin digit0<=ONE; digit1<=SEVEN; digit2<=SIX; digit3<=SEVEN; end
      16'd7672: begin digit0<=TWO; digit1<=SEVEN; digit2<=SIX; digit3<=SEVEN; end
      16'd7673: begin digit0<=THREE; digit1<=SEVEN; digit2<=SIX; digit3<=SEVEN; end
      16'd7674: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SIX; digit3<=SEVEN; end
      16'd7675: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SIX; digit3<=SEVEN; end
      16'd7676: begin digit0<=SIX; digit1<=SEVEN; digit2<=SIX; digit3<=SEVEN; end
      16'd7677: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SIX; digit3<=SEVEN; end
      16'd7678: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SIX; digit3<=SEVEN; end
      16'd7679: begin digit0<=NINE; digit1<=SEVEN; digit2<=SIX; digit3<=SEVEN; end
      16'd7680: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=SEVEN; end
      16'd7681: begin digit0<=ONE; digit1<=EIGHT; digit2<=SIX; digit3<=SEVEN; end
      16'd7682: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=SEVEN; end
      16'd7683: begin digit0<=THREE; digit1<=EIGHT; digit2<=SIX; digit3<=SEVEN; end
      16'd7684: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SIX; digit3<=SEVEN; end
      16'd7685: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SIX; digit3<=SEVEN; end
      16'd7686: begin digit0<=SIX; digit1<=EIGHT; digit2<=SIX; digit3<=SEVEN; end
      16'd7687: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SIX; digit3<=SEVEN; end
      16'd7688: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SIX; digit3<=SEVEN; end
      16'd7689: begin digit0<=NINE; digit1<=EIGHT; digit2<=SIX; digit3<=SEVEN; end
      16'd7690: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=SEVEN; end
      16'd7691: begin digit0<=ONE; digit1<=NINE; digit2<=SIX; digit3<=SEVEN; end
      16'd7692: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=SEVEN; end
      16'd7693: begin digit0<=THREE; digit1<=NINE; digit2<=SIX; digit3<=SEVEN; end
      16'd7694: begin digit0<=FOUR; digit1<=NINE; digit2<=SIX; digit3<=SEVEN; end
      16'd7695: begin digit0<=FIVE; digit1<=NINE; digit2<=SIX; digit3<=SEVEN; end
      16'd7696: begin digit0<=SIX; digit1<=NINE; digit2<=SIX; digit3<=SEVEN; end
      16'd7697: begin digit0<=SEVEN; digit1<=NINE; digit2<=SIX; digit3<=SEVEN; end
      16'd7698: begin digit0<=EIGHT; digit1<=NINE; digit2<=SIX; digit3<=SEVEN; end
      16'd7699: begin digit0<=NINE; digit1<=NINE; digit2<=SIX; digit3<=SEVEN; end
	  16'd7700: begin digit0<=ZERO; digit1<=ZERO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7701: begin digit0<=ONE; digit1<=ZERO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7702: begin digit0<=TWO; digit1<=ZERO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7703: begin digit0<=THREE; digit1<=ZERO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7704: begin digit0<=FOUR; digit1<=ZERO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7705: begin digit0<=FIVE; digit1<=ZERO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7706: begin digit0<=SIX; digit1<=ZERO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7707: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7708: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7709: begin digit0<=NINE; digit1<=ZERO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7710: begin digit0<=ZERO; digit1<=ONE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7711: begin digit0<=ONE; digit1<=ONE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7712: begin digit0<=TWO; digit1<=ONE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7713: begin digit0<=THREE; digit1<=ONE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7714: begin digit0<=FOUR; digit1<=ONE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7715: begin digit0<=FIVE; digit1<=ONE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7716: begin digit0<=SIX; digit1<=ONE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7717: begin digit0<=SEVEN; digit1<=ONE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7718: begin digit0<=EIGHT; digit1<=ONE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7719: begin digit0<=NINE; digit1<=ONE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7720: begin digit0<=ZERO; digit1<=TWO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7721: begin digit0<=ONE; digit1<=TWO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7722: begin digit0<=TWO; digit1<=TWO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7723: begin digit0<=THREE; digit1<=TWO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7724: begin digit0<=FOUR; digit1<=TWO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7725: begin digit0<=FIVE; digit1<=TWO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7726: begin digit0<=SIX; digit1<=TWO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7727: begin digit0<=SEVEN; digit1<=TWO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7728: begin digit0<=EIGHT; digit1<=TWO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7729: begin digit0<=NINE; digit1<=TWO; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7730: begin digit0<=ZERO; digit1<=THREE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7731: begin digit0<=ONE; digit1<=THREE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7732: begin digit0<=TWO; digit1<=THREE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7733: begin digit0<=THREE; digit1<=THREE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7734: begin digit0<=FOUR; digit1<=THREE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7735: begin digit0<=FIVE; digit1<=THREE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7736: begin digit0<=SIX; digit1<=THREE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7737: begin digit0<=SEVEN; digit1<=THREE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7738: begin digit0<=EIGHT; digit1<=THREE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7739: begin digit0<=NINE; digit1<=THREE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7740: begin digit0<=ZERO; digit1<=FOUR; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7741: begin digit0<=ONE; digit1<=FOUR; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7742: begin digit0<=TWO; digit1<=FOUR; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7743: begin digit0<=THREE; digit1<=FOUR; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7744: begin digit0<=FOUR; digit1<=FOUR; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7745: begin digit0<=FIVE; digit1<=FOUR; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7746: begin digit0<=SIX; digit1<=FOUR; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7747: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7748: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7749: begin digit0<=NINE; digit1<=FOUR; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7750: begin digit0<=ZERO; digit1<=FIVE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7751: begin digit0<=ONE; digit1<=FIVE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7752: begin digit0<=TWO; digit1<=FIVE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7753: begin digit0<=THREE; digit1<=FIVE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7754: begin digit0<=FOUR; digit1<=FIVE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7755: begin digit0<=FIVE; digit1<=FIVE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7756: begin digit0<=SIX; digit1<=FIVE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7757: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7758: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7759: begin digit0<=NINE; digit1<=FIVE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7760: begin digit0<=ZERO; digit1<=SIX; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7761: begin digit0<=ONE; digit1<=SIX; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7762: begin digit0<=TWO; digit1<=SIX; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7763: begin digit0<=THREE; digit1<=SIX; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7764: begin digit0<=FOUR; digit1<=SIX; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7765: begin digit0<=FIVE; digit1<=SIX; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7766: begin digit0<=SIX; digit1<=SIX; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7767: begin digit0<=SEVEN; digit1<=SIX; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7768: begin digit0<=EIGHT; digit1<=SIX; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7769: begin digit0<=NINE; digit1<=SIX; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7770: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7771: begin digit0<=ONE; digit1<=SEVEN; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7772: begin digit0<=TWO; digit1<=SEVEN; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7773: begin digit0<=THREE; digit1<=SEVEN; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7774: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7775: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7776: begin digit0<=SIX; digit1<=SEVEN; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7777: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7778: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7779: begin digit0<=NINE; digit1<=SEVEN; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7780: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7781: begin digit0<=ONE; digit1<=EIGHT; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7782: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7783: begin digit0<=THREE; digit1<=EIGHT; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7784: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7785: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7786: begin digit0<=SIX; digit1<=EIGHT; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7787: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7788: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7789: begin digit0<=NINE; digit1<=EIGHT; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7790: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7791: begin digit0<=ONE; digit1<=NINE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7792: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7793: begin digit0<=THREE; digit1<=NINE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7794: begin digit0<=FOUR; digit1<=NINE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7795: begin digit0<=FIVE; digit1<=NINE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7796: begin digit0<=SIX; digit1<=NINE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7797: begin digit0<=SEVEN; digit1<=NINE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7798: begin digit0<=EIGHT; digit1<=NINE; digit2<=SEVEN; digit3<=SEVEN; end
      16'd7799: begin digit0<=NINE; digit1<=NINE; digit2<=SEVEN; digit3<=SEVEN; end
	  16'd7800: begin digit0<=ZERO; digit1<=ZERO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7801: begin digit0<=ONE; digit1<=ZERO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7802: begin digit0<=TWO; digit1<=ZERO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7803: begin digit0<=THREE; digit1<=ZERO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7804: begin digit0<=FOUR; digit1<=ZERO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7805: begin digit0<=FIVE; digit1<=ZERO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7806: begin digit0<=SIX; digit1<=ZERO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7807: begin digit0<=SEVEN; digit1<=ZERO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7808: begin digit0<=EIGHT; digit1<=ZERO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7809: begin digit0<=NINE; digit1<=ZERO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7810: begin digit0<=ZERO; digit1<=ONE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7811: begin digit0<=ONE; digit1<=ONE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7812: begin digit0<=TWO; digit1<=ONE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7813: begin digit0<=THREE; digit1<=ONE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7814: begin digit0<=FOUR; digit1<=ONE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7815: begin digit0<=FIVE; digit1<=ONE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7816: begin digit0<=SIX; digit1<=ONE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7817: begin digit0<=SEVEN; digit1<=ONE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7818: begin digit0<=EIGHT; digit1<=ONE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7819: begin digit0<=NINE; digit1<=ONE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7820: begin digit0<=ZERO; digit1<=TWO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7821: begin digit0<=ONE; digit1<=TWO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7822: begin digit0<=TWO; digit1<=TWO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7823: begin digit0<=THREE; digit1<=TWO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7824: begin digit0<=FOUR; digit1<=TWO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7825: begin digit0<=FIVE; digit1<=TWO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7826: begin digit0<=SIX; digit1<=TWO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7827: begin digit0<=SEVEN; digit1<=TWO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7828: begin digit0<=EIGHT; digit1<=TWO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7829: begin digit0<=NINE; digit1<=TWO; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7830: begin digit0<=ZERO; digit1<=THREE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7831: begin digit0<=ONE; digit1<=THREE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7832: begin digit0<=TWO; digit1<=THREE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7833: begin digit0<=THREE; digit1<=THREE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7834: begin digit0<=FOUR; digit1<=THREE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7835: begin digit0<=FIVE; digit1<=THREE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7836: begin digit0<=SIX; digit1<=THREE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7837: begin digit0<=SEVEN; digit1<=THREE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7838: begin digit0<=EIGHT; digit1<=THREE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7839: begin digit0<=NINE; digit1<=THREE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7840: begin digit0<=ZERO; digit1<=FOUR; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7841: begin digit0<=ONE; digit1<=FOUR; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7842: begin digit0<=TWO; digit1<=FOUR; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7843: begin digit0<=THREE; digit1<=FOUR; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7844: begin digit0<=FOUR; digit1<=FOUR; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7845: begin digit0<=FIVE; digit1<=FOUR; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7846: begin digit0<=SIX; digit1<=FOUR; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7847: begin digit0<=SEVEN; digit1<=FOUR; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7848: begin digit0<=EIGHT; digit1<=FOUR; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7849: begin digit0<=NINE; digit1<=FOUR; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7850: begin digit0<=ZERO; digit1<=FIVE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7851: begin digit0<=ONE; digit1<=FIVE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7852: begin digit0<=TWO; digit1<=FIVE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7853: begin digit0<=THREE; digit1<=FIVE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7854: begin digit0<=FOUR; digit1<=FIVE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7855: begin digit0<=FIVE; digit1<=FIVE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7856: begin digit0<=SIX; digit1<=FIVE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7857: begin digit0<=SEVEN; digit1<=FIVE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7858: begin digit0<=EIGHT; digit1<=FIVE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7859: begin digit0<=NINE; digit1<=FIVE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7860: begin digit0<=ZERO; digit1<=SIX; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7861: begin digit0<=ONE; digit1<=SIX; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7862: begin digit0<=TWO; digit1<=SIX; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7863: begin digit0<=THREE; digit1<=SIX; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7864: begin digit0<=FOUR; digit1<=SIX; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7865: begin digit0<=FIVE; digit1<=SIX; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7866: begin digit0<=SIX; digit1<=SIX; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7867: begin digit0<=SEVEN; digit1<=SIX; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7868: begin digit0<=EIGHT; digit1<=SIX; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7869: begin digit0<=NINE; digit1<=SIX; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7870: begin digit0<=ZERO; digit1<=SEVEN; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7871: begin digit0<=ONE; digit1<=SEVEN; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7872: begin digit0<=TWO; digit1<=SEVEN; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7873: begin digit0<=THREE; digit1<=SEVEN; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7874: begin digit0<=FOUR; digit1<=SEVEN; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7875: begin digit0<=FIVE; digit1<=SEVEN; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7876: begin digit0<=SIX; digit1<=SEVEN; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7877: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7878: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7879: begin digit0<=NINE; digit1<=SEVEN; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7880: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7881: begin digit0<=ONE; digit1<=EIGHT; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7882: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7883: begin digit0<=THREE; digit1<=EIGHT; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7884: begin digit0<=FOUR; digit1<=EIGHT; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7885: begin digit0<=FIVE; digit1<=EIGHT; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7886: begin digit0<=SIX; digit1<=EIGHT; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7887: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7888: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7889: begin digit0<=NINE; digit1<=EIGHT; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7890: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7891: begin digit0<=ONE; digit1<=NINE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7892: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7893: begin digit0<=THREE; digit1<=NINE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7894: begin digit0<=FOUR; digit1<=NINE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7895: begin digit0<=FIVE; digit1<=NINE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7896: begin digit0<=SIX; digit1<=NINE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7897: begin digit0<=SEVEN; digit1<=NINE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7898: begin digit0<=EIGHT; digit1<=NINE; digit2<=EIGHT; digit3<=SEVEN; end
      16'd7899: begin digit0<=NINE; digit1<=NINE; digit2<=EIGHT; digit3<=SEVEN; end
	  16'd7900: begin digit0<=ZERO; digit1<=ZERO; digit2<=NINE; digit3<=SEVEN; end
      16'd7901: begin digit0<=ONE; digit1<=ZERO; digit2<=NINE; digit3<=SEVEN; end
      16'd7902: begin digit0<=TWO; digit1<=ZERO; digit2<=NINE; digit3<=SEVEN; end
      16'd7903: begin digit0<=THREE; digit1<=ZERO; digit2<=NINE; digit3<=SEVEN; end
      16'd7904: begin digit0<=FOUR; digit1<=ZERO; digit2<=NINE; digit3<=SEVEN; end
      16'd7905: begin digit0<=FIVE; digit1<=ZERO; digit2<=NINE; digit3<=SEVEN; end
      16'd7906: begin digit0<=SIX; digit1<=ZERO; digit2<=NINE; digit3<=SEVEN; end
      16'd7907: begin digit0<=SEVEN; digit1<=ZERO; digit2<=NINE; digit3<=SEVEN; end
      16'd7908: begin digit0<=EIGHT; digit1<=ZERO; digit2<=NINE; digit3<=SEVEN; end
      16'd7909: begin digit0<=NINE; digit1<=ZERO; digit2<=NINE; digit3<=SEVEN; end
      16'd7910: begin digit0<=ZERO; digit1<=ONE; digit2<=NINE; digit3<=SEVEN; end
      16'd7911: begin digit0<=ONE; digit1<=ONE; digit2<=NINE; digit3<=SEVEN; end
      16'd7912: begin digit0<=TWO; digit1<=ONE; digit2<=NINE; digit3<=SEVEN; end
      16'd7913: begin digit0<=THREE; digit1<=ONE; digit2<=NINE; digit3<=SEVEN; end
      16'd7914: begin digit0<=FOUR; digit1<=ONE; digit2<=NINE; digit3<=SEVEN; end
      16'd7915: begin digit0<=FIVE; digit1<=ONE; digit2<=NINE; digit3<=SEVEN; end
      16'd7916: begin digit0<=SIX; digit1<=ONE; digit2<=NINE; digit3<=SEVEN; end
      16'd7917: begin digit0<=SEVEN; digit1<=ONE; digit2<=NINE; digit3<=SEVEN; end
      16'd7918: begin digit0<=EIGHT; digit1<=ONE; digit2<=NINE; digit3<=SEVEN; end
      16'd7919: begin digit0<=NINE; digit1<=ONE; digit2<=NINE; digit3<=SEVEN; end
      16'd7920: begin digit0<=ZERO; digit1<=TWO; digit2<=NINE; digit3<=SEVEN; end
      16'd7921: begin digit0<=ONE; digit1<=TWO; digit2<=NINE; digit3<=SEVEN; end
      16'd7922: begin digit0<=TWO; digit1<=TWO; digit2<=NINE; digit3<=SEVEN; end
      16'd7923: begin digit0<=THREE; digit1<=TWO; digit2<=NINE; digit3<=SEVEN; end
      16'd7924: begin digit0<=FOUR; digit1<=TWO; digit2<=NINE; digit3<=SEVEN; end
      16'd7925: begin digit0<=FIVE; digit1<=TWO; digit2<=NINE; digit3<=SEVEN; end
      16'd7926: begin digit0<=SIX; digit1<=TWO; digit2<=NINE; digit3<=SEVEN; end
      16'd7927: begin digit0<=SEVEN; digit1<=TWO; digit2<=NINE; digit3<=SEVEN; end
      16'd7928: begin digit0<=EIGHT; digit1<=TWO; digit2<=NINE; digit3<=SEVEN; end
      16'd7929: begin digit0<=NINE; digit1<=TWO; digit2<=NINE; digit3<=SEVEN; end
      16'd7930: begin digit0<=ZERO; digit1<=THREE; digit2<=NINE; digit3<=SEVEN; end
      16'd7931: begin digit0<=ONE; digit1<=THREE; digit2<=NINE; digit3<=SEVEN; end
      16'd7932: begin digit0<=TWO; digit1<=THREE; digit2<=NINE; digit3<=SEVEN; end
      16'd7933: begin digit0<=THREE; digit1<=THREE; digit2<=NINE; digit3<=SEVEN; end
      16'd7934: begin digit0<=FOUR; digit1<=THREE; digit2<=NINE; digit3<=SEVEN; end
      16'd7935: begin digit0<=FIVE; digit1<=THREE; digit2<=NINE; digit3<=SEVEN; end
      16'd7936: begin digit0<=SIX; digit1<=THREE; digit2<=NINE; digit3<=SEVEN; end
      16'd7937: begin digit0<=SEVEN; digit1<=THREE; digit2<=NINE; digit3<=SEVEN; end
      16'd7938: begin digit0<=EIGHT; digit1<=THREE; digit2<=NINE; digit3<=SEVEN; end
      16'd7939: begin digit0<=NINE; digit1<=THREE; digit2<=NINE; digit3<=SEVEN; end
      16'd7940: begin digit0<=ZERO; digit1<=FOUR; digit2<=NINE; digit3<=SEVEN; end
      16'd7941: begin digit0<=ONE; digit1<=FOUR; digit2<=NINE; digit3<=SEVEN; end
      16'd7942: begin digit0<=TWO; digit1<=FOUR; digit2<=NINE; digit3<=SEVEN; end
      16'd7943: begin digit0<=THREE; digit1<=FOUR; digit2<=NINE; digit3<=SEVEN; end
      16'd7944: begin digit0<=FOUR; digit1<=FOUR; digit2<=NINE; digit3<=SEVEN; end
      16'd7945: begin digit0<=FIVE; digit1<=FOUR; digit2<=NINE; digit3<=SEVEN; end
      16'd7946: begin digit0<=SIX; digit1<=FOUR; digit2<=NINE; digit3<=SEVEN; end
      16'd7947: begin digit0<=SEVEN; digit1<=FOUR; digit2<=NINE; digit3<=SEVEN; end
      16'd7948: begin digit0<=EIGHT; digit1<=FOUR; digit2<=NINE; digit3<=SEVEN; end
      16'd7949: begin digit0<=NINE; digit1<=FOUR; digit2<=NINE; digit3<=SEVEN; end
      16'd7950: begin digit0<=ZERO; digit1<=FIVE; digit2<=NINE; digit3<=SEVEN; end
      16'd7951: begin digit0<=ONE; digit1<=FIVE; digit2<=NINE; digit3<=SEVEN; end
      16'd7952: begin digit0<=TWO; digit1<=FIVE; digit2<=NINE; digit3<=SEVEN; end
      16'd7953: begin digit0<=THREE; digit1<=FIVE; digit2<=NINE; digit3<=SEVEN; end
      16'd7954: begin digit0<=FOUR; digit1<=FIVE; digit2<=NINE; digit3<=SEVEN; end
      16'd7955: begin digit0<=FIVE; digit1<=FIVE; digit2<=NINE; digit3<=SEVEN; end
      16'd7956: begin digit0<=SIX; digit1<=FIVE; digit2<=NINE; digit3<=SEVEN; end
      16'd7957: begin digit0<=SEVEN; digit1<=FIVE; digit2<=NINE; digit3<=SEVEN; end
      16'd7958: begin digit0<=EIGHT; digit1<=FIVE; digit2<=NINE; digit3<=SEVEN; end
      16'd7959: begin digit0<=NINE; digit1<=FIVE; digit2<=NINE; digit3<=SEVEN; end
      16'd7960: begin digit0<=ZERO; digit1<=SIX; digit2<=NINE; digit3<=SEVEN; end
      16'd7961: begin digit0<=ONE; digit1<=SIX; digit2<=NINE; digit3<=SEVEN; end
      16'd7962: begin digit0<=TWO; digit1<=SIX; digit2<=NINE; digit3<=SEVEN; end
      16'd7963: begin digit0<=THREE; digit1<=SIX; digit2<=NINE; digit3<=SEVEN; end
      16'd7964: begin digit0<=FOUR; digit1<=SIX; digit2<=NINE; digit3<=SEVEN; end
      16'd7965: begin digit0<=FIVE; digit1<=SIX; digit2<=NINE; digit3<=SEVEN; end
      16'd7966: begin digit0<=SIX; digit1<=SIX; digit2<=NINE; digit3<=SEVEN; end
      16'd7967: begin digit0<=SEVEN; digit1<=SIX; digit2<=NINE; digit3<=SEVEN; end
      16'd7968: begin digit0<=EIGHT; digit1<=SIX; digit2<=NINE; digit3<=SEVEN; end
      16'd7969: begin digit0<=NINE; digit1<=SIX; digit2<=NINE; digit3<=SEVEN; end
      16'd7970: begin digit0<=ZERO; digit1<=SEVEN; digit2<=NINE; digit3<=SEVEN; end
      16'd7971: begin digit0<=ONE; digit1<=SEVEN; digit2<=NINE; digit3<=SEVEN; end
      16'd7972: begin digit0<=TWO; digit1<=SEVEN; digit2<=NINE; digit3<=SEVEN; end
      16'd7973: begin digit0<=THREE; digit1<=SEVEN; digit2<=NINE; digit3<=SEVEN; end
      16'd7974: begin digit0<=FOUR; digit1<=SEVEN; digit2<=NINE; digit3<=SEVEN; end
      16'd7975: begin digit0<=FIVE; digit1<=SEVEN; digit2<=NINE; digit3<=SEVEN; end
      16'd7976: begin digit0<=SIX; digit1<=SEVEN; digit2<=NINE; digit3<=SEVEN; end
      16'd7977: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=NINE; digit3<=SEVEN; end
      16'd7978: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=NINE; digit3<=SEVEN; end
      16'd7979: begin digit0<=NINE; digit1<=SEVEN; digit2<=NINE; digit3<=SEVEN; end
      16'd7980: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=SEVEN; end
      16'd7981: begin digit0<=ONE; digit1<=EIGHT; digit2<=NINE; digit3<=SEVEN; end
      16'd7982: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=SEVEN; end
      16'd7983: begin digit0<=THREE; digit1<=EIGHT; digit2<=NINE; digit3<=SEVEN; end
      16'd7984: begin digit0<=FOUR; digit1<=EIGHT; digit2<=NINE; digit3<=SEVEN; end
      16'd7985: begin digit0<=FIVE; digit1<=EIGHT; digit2<=NINE; digit3<=SEVEN; end
      16'd7986: begin digit0<=SIX; digit1<=EIGHT; digit2<=NINE; digit3<=SEVEN; end
      16'd7987: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=NINE; digit3<=SEVEN; end
      16'd7988: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=NINE; digit3<=SEVEN; end
      16'd7989: begin digit0<=NINE; digit1<=EIGHT; digit2<=NINE; digit3<=SEVEN; end
      16'd7990: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=SEVEN; end
      16'd7991: begin digit0<=ONE; digit1<=NINE; digit2<=NINE; digit3<=SEVEN; end
      16'd7992: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=SEVEN; end
      16'd7993: begin digit0<=THREE; digit1<=NINE; digit2<=NINE; digit3<=SEVEN; end
      16'd7994: begin digit0<=FOUR; digit1<=NINE; digit2<=NINE; digit3<=SEVEN; end
      16'd7995: begin digit0<=FIVE; digit1<=NINE; digit2<=NINE; digit3<=SEVEN; end
      16'd7996: begin digit0<=SIX; digit1<=NINE; digit2<=NINE; digit3<=SEVEN; end
      16'd7997: begin digit0<=SEVEN; digit1<=NINE; digit2<=NINE; digit3<=SEVEN; end
      16'd7998: begin digit0<=EIGHT; digit1<=NINE; digit2<=NINE; digit3<=SEVEN; end
      16'd7999: begin digit0<=NINE; digit1<=NINE; digit2<=NINE; digit3<=SEVEN; end
	  16'd8000: begin digit0<=ZERO; digit1<=ZERO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8001: begin digit0<=ONE; digit1<=ZERO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8002: begin digit0<=TWO; digit1<=ZERO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8003: begin digit0<=THREE; digit1<=ZERO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8004: begin digit0<=FOUR; digit1<=ZERO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8005: begin digit0<=FIVE; digit1<=ZERO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8006: begin digit0<=SIX; digit1<=ZERO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8007: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8008: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8009: begin digit0<=NINE; digit1<=ZERO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8010: begin digit0<=ZERO; digit1<=ONE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8011: begin digit0<=ONE; digit1<=ONE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8012: begin digit0<=TWO; digit1<=ONE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8013: begin digit0<=THREE; digit1<=ONE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8014: begin digit0<=FOUR; digit1<=ONE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8015: begin digit0<=FIVE; digit1<=ONE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8016: begin digit0<=SIX; digit1<=ONE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8017: begin digit0<=SEVEN; digit1<=ONE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8018: begin digit0<=EIGHT; digit1<=ONE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8019: begin digit0<=NINE; digit1<=ONE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8020: begin digit0<=ZERO; digit1<=TWO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8021: begin digit0<=ONE; digit1<=TWO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8022: begin digit0<=TWO; digit1<=TWO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8023: begin digit0<=THREE; digit1<=TWO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8024: begin digit0<=FOUR; digit1<=TWO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8025: begin digit0<=FIVE; digit1<=TWO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8026: begin digit0<=SIX; digit1<=TWO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8027: begin digit0<=SEVEN; digit1<=TWO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8028: begin digit0<=EIGHT; digit1<=TWO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8029: begin digit0<=NINE; digit1<=TWO; digit2<=ZERO; digit3<=EIGHT; end
      16'd8030: begin digit0<=ZERO; digit1<=THREE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8031: begin digit0<=ONE; digit1<=THREE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8032: begin digit0<=TWO; digit1<=THREE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8033: begin digit0<=THREE; digit1<=THREE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8034: begin digit0<=FOUR; digit1<=THREE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8035: begin digit0<=FIVE; digit1<=THREE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8036: begin digit0<=SIX; digit1<=THREE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8037: begin digit0<=SEVEN; digit1<=THREE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8038: begin digit0<=EIGHT; digit1<=THREE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8039: begin digit0<=NINE; digit1<=THREE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8040: begin digit0<=ZERO; digit1<=FOUR; digit2<=ZERO; digit3<=EIGHT; end
      16'd8041: begin digit0<=ONE; digit1<=FOUR; digit2<=ZERO; digit3<=EIGHT; end
      16'd8042: begin digit0<=TWO; digit1<=FOUR; digit2<=ZERO; digit3<=EIGHT; end
      16'd8043: begin digit0<=THREE; digit1<=FOUR; digit2<=ZERO; digit3<=EIGHT; end
      16'd8044: begin digit0<=FOUR; digit1<=FOUR; digit2<=ZERO; digit3<=EIGHT; end
      16'd8045: begin digit0<=FIVE; digit1<=FOUR; digit2<=ZERO; digit3<=EIGHT; end
      16'd8046: begin digit0<=SIX; digit1<=FOUR; digit2<=ZERO; digit3<=EIGHT; end
      16'd8047: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ZERO; digit3<=EIGHT; end
      16'd8048: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ZERO; digit3<=EIGHT; end
      16'd8049: begin digit0<=NINE; digit1<=FOUR; digit2<=ZERO; digit3<=EIGHT; end
      16'd8050: begin digit0<=ZERO; digit1<=FIVE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8051: begin digit0<=ONE; digit1<=FIVE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8052: begin digit0<=TWO; digit1<=FIVE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8053: begin digit0<=THREE; digit1<=FIVE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8054: begin digit0<=FOUR; digit1<=FIVE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8055: begin digit0<=FIVE; digit1<=FIVE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8056: begin digit0<=SIX; digit1<=FIVE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8057: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8058: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8059: begin digit0<=NINE; digit1<=FIVE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8060: begin digit0<=ZERO; digit1<=SIX; digit2<=ZERO; digit3<=EIGHT; end
      16'd8061: begin digit0<=ONE; digit1<=SIX; digit2<=ZERO; digit3<=EIGHT; end
      16'd8062: begin digit0<=TWO; digit1<=SIX; digit2<=ZERO; digit3<=EIGHT; end
      16'd8063: begin digit0<=THREE; digit1<=SIX; digit2<=ZERO; digit3<=EIGHT; end
      16'd8064: begin digit0<=FOUR; digit1<=SIX; digit2<=ZERO; digit3<=EIGHT; end
      16'd8065: begin digit0<=FIVE; digit1<=SIX; digit2<=ZERO; digit3<=EIGHT; end
      16'd8066: begin digit0<=SIX; digit1<=SIX; digit2<=ZERO; digit3<=EIGHT; end
      16'd8067: begin digit0<=SEVEN; digit1<=SIX; digit2<=ZERO; digit3<=EIGHT; end
      16'd8068: begin digit0<=EIGHT; digit1<=SIX; digit2<=ZERO; digit3<=EIGHT; end
      16'd8069: begin digit0<=NINE; digit1<=SIX; digit2<=ZERO; digit3<=EIGHT; end
      16'd8070: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ZERO; digit3<=EIGHT; end
      16'd8071: begin digit0<=ONE; digit1<=SEVEN; digit2<=ZERO; digit3<=EIGHT; end
      16'd8072: begin digit0<=TWO; digit1<=SEVEN; digit2<=ZERO; digit3<=EIGHT; end
      16'd8073: begin digit0<=THREE; digit1<=SEVEN; digit2<=ZERO; digit3<=EIGHT; end
      16'd8074: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ZERO; digit3<=EIGHT; end
      16'd8075: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ZERO; digit3<=EIGHT; end
      16'd8076: begin digit0<=SIX; digit1<=SEVEN; digit2<=ZERO; digit3<=EIGHT; end
      16'd8077: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ZERO; digit3<=EIGHT; end
      16'd8078: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ZERO; digit3<=EIGHT; end
      16'd8079: begin digit0<=NINE; digit1<=SEVEN; digit2<=ZERO; digit3<=EIGHT; end
      16'd8080: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ZERO; digit3<=EIGHT; end
      16'd8081: begin digit0<=ONE; digit1<=EIGHT; digit2<=ZERO; digit3<=EIGHT; end
      16'd8082: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ZERO; digit3<=EIGHT; end
      16'd8083: begin digit0<=THREE; digit1<=EIGHT; digit2<=ZERO; digit3<=EIGHT; end
      16'd8084: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ZERO; digit3<=EIGHT; end
      16'd8085: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ZERO; digit3<=EIGHT; end
      16'd8086: begin digit0<=SIX; digit1<=EIGHT; digit2<=ZERO; digit3<=EIGHT; end
      16'd8087: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ZERO; digit3<=EIGHT; end
      16'd8088: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ZERO; digit3<=EIGHT; end
      16'd8089: begin digit0<=NINE; digit1<=EIGHT; digit2<=ZERO; digit3<=EIGHT; end
      16'd8090: begin digit0<=ZERO; digit1<=NINE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8091: begin digit0<=ONE; digit1<=NINE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8092: begin digit0<=ZERO; digit1<=NINE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8093: begin digit0<=THREE; digit1<=NINE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8094: begin digit0<=FOUR; digit1<=NINE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8095: begin digit0<=FIVE; digit1<=NINE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8096: begin digit0<=SIX; digit1<=NINE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8097: begin digit0<=SEVEN; digit1<=NINE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8098: begin digit0<=EIGHT; digit1<=NINE; digit2<=ZERO; digit3<=EIGHT; end
      16'd8099: begin digit0<=NINE; digit1<=NINE; digit2<=ZERO; digit3<=EIGHT; end
	  16'd8100: begin digit0<=ZERO; digit1<=ZERO; digit2<=ONE; digit3<=EIGHT; end
      16'd8101: begin digit0<=ONE; digit1<=ZERO; digit2<=ONE; digit3<=EIGHT; end
      16'd8102: begin digit0<=TWO; digit1<=ZERO; digit2<=ONE; digit3<=EIGHT; end
      16'd8103: begin digit0<=THREE; digit1<=ZERO; digit2<=ONE; digit3<=EIGHT; end
      16'd8104: begin digit0<=FOUR; digit1<=ZERO; digit2<=ONE; digit3<=EIGHT; end
      16'd8105: begin digit0<=FIVE; digit1<=ZERO; digit2<=ONE; digit3<=EIGHT; end
      16'd8106: begin digit0<=SIX; digit1<=ZERO; digit2<=ONE; digit3<=EIGHT; end
      16'd8107: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ONE; digit3<=EIGHT; end
      16'd8108: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ONE; digit3<=EIGHT; end
      16'd8109: begin digit0<=NINE; digit1<=ZERO; digit2<=ONE; digit3<=EIGHT; end
      16'd8110: begin digit0<=ZERO; digit1<=ONE; digit2<=ONE; digit3<=EIGHT; end
      16'd8111: begin digit0<=ONE; digit1<=ONE; digit2<=ONE; digit3<=EIGHT; end
      16'd8112: begin digit0<=TWO; digit1<=ONE; digit2<=ONE; digit3<=EIGHT; end
      16'd8113: begin digit0<=THREE; digit1<=ONE; digit2<=ONE; digit3<=EIGHT; end
      16'd8114: begin digit0<=FOUR; digit1<=ONE; digit2<=ONE; digit3<=EIGHT; end
      16'd8115: begin digit0<=FIVE; digit1<=ONE; digit2<=ONE; digit3<=EIGHT; end
      16'd8116: begin digit0<=SIX; digit1<=ONE; digit2<=ONE; digit3<=EIGHT; end
      16'd8117: begin digit0<=SEVEN; digit1<=ONE; digit2<=ONE; digit3<=EIGHT; end
      16'd8118: begin digit0<=EIGHT; digit1<=ONE; digit2<=ONE; digit3<=EIGHT; end
      16'd8119: begin digit0<=NINE; digit1<=ONE; digit2<=ONE; digit3<=EIGHT; end
      16'd8120: begin digit0<=ZERO; digit1<=TWO; digit2<=ONE; digit3<=EIGHT; end
      16'd8121: begin digit0<=ONE; digit1<=TWO; digit2<=ONE; digit3<=EIGHT; end
      16'd8122: begin digit0<=TWO; digit1<=TWO; digit2<=ONE; digit3<=EIGHT; end
      16'd8123: begin digit0<=THREE; digit1<=TWO; digit2<=ONE; digit3<=EIGHT; end
      16'd8124: begin digit0<=FOUR; digit1<=TWO; digit2<=ONE; digit3<=EIGHT; end
      16'd8125: begin digit0<=FIVE; digit1<=TWO; digit2<=ONE; digit3<=EIGHT; end
      16'd8126: begin digit0<=SIX; digit1<=TWO; digit2<=ONE; digit3<=EIGHT; end
      16'd8127: begin digit0<=SEVEN; digit1<=TWO; digit2<=ONE; digit3<=EIGHT; end
      16'd8128: begin digit0<=EIGHT; digit1<=TWO; digit2<=ONE; digit3<=EIGHT; end
      16'd8129: begin digit0<=NINE; digit1<=TWO; digit2<=ONE; digit3<=EIGHT; end
      16'd8130: begin digit0<=ZERO; digit1<=THREE; digit2<=ONE; digit3<=EIGHT; end
      16'd8131: begin digit0<=ONE; digit1<=THREE; digit2<=ONE; digit3<=EIGHT; end
      16'd8132: begin digit0<=TWO; digit1<=THREE; digit2<=ONE; digit3<=EIGHT; end
      16'd8133: begin digit0<=THREE; digit1<=THREE; digit2<=ONE; digit3<=EIGHT; end
      16'd8134: begin digit0<=FOUR; digit1<=THREE; digit2<=ONE; digit3<=EIGHT; end
      16'd8135: begin digit0<=FIVE; digit1<=THREE; digit2<=ONE; digit3<=EIGHT; end
      16'd8136: begin digit0<=SIX; digit1<=THREE; digit2<=ONE; digit3<=EIGHT; end
      16'd8137: begin digit0<=SEVEN; digit1<=THREE; digit2<=ONE; digit3<=EIGHT; end
      16'd8138: begin digit0<=EIGHT; digit1<=THREE; digit2<=ONE; digit3<=EIGHT; end
      16'd8139: begin digit0<=NINE; digit1<=THREE; digit2<=ONE; digit3<=EIGHT; end
      16'd8140: begin digit0<=ZERO; digit1<=FOUR; digit2<=ONE; digit3<=EIGHT; end
      16'd8141: begin digit0<=ONE; digit1<=FOUR; digit2<=ONE; digit3<=EIGHT; end
      16'd8142: begin digit0<=TWO; digit1<=FOUR; digit2<=ONE; digit3<=EIGHT; end
      16'd8143: begin digit0<=THREE; digit1<=FOUR; digit2<=ONE; digit3<=EIGHT; end
      16'd8144: begin digit0<=FOUR; digit1<=FOUR; digit2<=ONE; digit3<=EIGHT; end
      16'd8145: begin digit0<=FIVE; digit1<=FOUR; digit2<=ONE; digit3<=EIGHT; end
      16'd8146: begin digit0<=SIX; digit1<=FOUR; digit2<=ONE; digit3<=EIGHT; end
      16'd8147: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ONE; digit3<=EIGHT; end
      16'd8148: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ONE; digit3<=EIGHT; end
      16'd8149: begin digit0<=NINE; digit1<=FOUR; digit2<=ONE; digit3<=EIGHT; end
      16'd8150: begin digit0<=ZERO; digit1<=FIVE; digit2<=ONE; digit3<=EIGHT; end
      16'd8151: begin digit0<=ONE; digit1<=FIVE; digit2<=ONE; digit3<=EIGHT; end
      16'd8152: begin digit0<=TWO; digit1<=FIVE; digit2<=ONE; digit3<=EIGHT; end
      16'd8153: begin digit0<=THREE; digit1<=FIVE; digit2<=ONE; digit3<=EIGHT; end
      16'd8154: begin digit0<=FOUR; digit1<=FIVE; digit2<=ONE; digit3<=EIGHT; end
      16'd8155: begin digit0<=FIVE; digit1<=FIVE; digit2<=ONE; digit3<=EIGHT; end
      16'd8156: begin digit0<=SIX; digit1<=FIVE; digit2<=ONE; digit3<=EIGHT; end
      16'd8157: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ONE; digit3<=EIGHT; end
      16'd8158: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ONE; digit3<=EIGHT; end
      16'd8159: begin digit0<=NINE; digit1<=FIVE; digit2<=ONE; digit3<=EIGHT; end
      16'd8160: begin digit0<=ZERO; digit1<=SIX; digit2<=ONE; digit3<=EIGHT; end
      16'd8161: begin digit0<=ONE; digit1<=SIX; digit2<=ONE; digit3<=EIGHT; end
      16'd8162: begin digit0<=TWO; digit1<=SIX; digit2<=ONE; digit3<=EIGHT; end
      16'd8163: begin digit0<=THREE; digit1<=SIX; digit2<=ONE; digit3<=EIGHT; end
      16'd8164: begin digit0<=FOUR; digit1<=SIX; digit2<=ONE; digit3<=EIGHT; end
      16'd8165: begin digit0<=FIVE; digit1<=SIX; digit2<=ONE; digit3<=EIGHT; end
      16'd8166: begin digit0<=SIX; digit1<=SIX; digit2<=ONE; digit3<=EIGHT; end
      16'd8167: begin digit0<=SEVEN; digit1<=SIX; digit2<=ONE; digit3<=EIGHT; end
      16'd8168: begin digit0<=EIGHT; digit1<=SIX; digit2<=ONE; digit3<=EIGHT; end
      16'd8169: begin digit0<=NINE; digit1<=SIX; digit2<=ONE; digit3<=EIGHT; end
      16'd8170: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ONE; digit3<=EIGHT; end
      16'd8171: begin digit0<=ONE; digit1<=SEVEN; digit2<=ONE; digit3<=EIGHT; end
      16'd8172: begin digit0<=TWO; digit1<=SEVEN; digit2<=ONE; digit3<=EIGHT; end
      16'd8173: begin digit0<=THREE; digit1<=SEVEN; digit2<=ONE; digit3<=EIGHT; end
      16'd8174: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ONE; digit3<=EIGHT; end
      16'd8175: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ONE; digit3<=EIGHT; end
      16'd8176: begin digit0<=SIX; digit1<=SEVEN; digit2<=ONE; digit3<=EIGHT; end
      16'd8177: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ONE; digit3<=EIGHT; end
      16'd8178: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ONE; digit3<=EIGHT; end
      16'd8179: begin digit0<=NINE; digit1<=SEVEN; digit2<=ONE; digit3<=EIGHT; end
      16'd8180: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=EIGHT; end
      16'd8181: begin digit0<=ONE; digit1<=EIGHT; digit2<=ONE; digit3<=EIGHT; end
      16'd8182: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=EIGHT; end
      16'd8183: begin digit0<=THREE; digit1<=EIGHT; digit2<=ONE; digit3<=EIGHT; end
      16'd8184: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ONE; digit3<=EIGHT; end
      16'd8185: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ONE; digit3<=EIGHT; end
      16'd8186: begin digit0<=SIX; digit1<=EIGHT; digit2<=ONE; digit3<=EIGHT; end
      16'd8187: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ONE; digit3<=EIGHT; end
      16'd8188: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ONE; digit3<=EIGHT; end
      16'd8189: begin digit0<=NINE; digit1<=EIGHT; digit2<=ONE; digit3<=EIGHT; end
      16'd8190: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=EIGHT; end
      16'd8191: begin digit0<=ONE; digit1<=NINE; digit2<=ONE; digit3<=EIGHT; end
      16'd8192: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=EIGHT; end
      16'd8193: begin digit0<=THREE; digit1<=NINE; digit2<=ONE; digit3<=EIGHT; end
      16'd8194: begin digit0<=FOUR; digit1<=NINE; digit2<=ONE; digit3<=EIGHT; end
      16'd8195: begin digit0<=FIVE; digit1<=NINE; digit2<=ONE; digit3<=EIGHT; end
      16'd8196: begin digit0<=SIX; digit1<=NINE; digit2<=ONE; digit3<=EIGHT; end
      16'd8197: begin digit0<=SEVEN; digit1<=NINE; digit2<=ONE; digit3<=EIGHT; end
      16'd8198: begin digit0<=EIGHT; digit1<=NINE; digit2<=ONE; digit3<=EIGHT; end
      16'd8199: begin digit0<=NINE; digit1<=NINE; digit2<=ONE; digit3<=EIGHT; end
	  16'd8200: begin digit0<=ZERO; digit1<=ZERO; digit2<=TWO; digit3<=EIGHT; end
      16'd8201: begin digit0<=ONE; digit1<=ZERO; digit2<=TWO; digit3<=EIGHT; end
      16'd8202: begin digit0<=TWO; digit1<=ZERO; digit2<=TWO; digit3<=EIGHT; end
      16'd8203: begin digit0<=THREE; digit1<=ZERO; digit2<=TWO; digit3<=EIGHT; end
      16'd8204: begin digit0<=FOUR; digit1<=ZERO; digit2<=TWO; digit3<=EIGHT; end
      16'd8205: begin digit0<=FIVE; digit1<=ZERO; digit2<=TWO; digit3<=EIGHT; end
      16'd8206: begin digit0<=SIX; digit1<=ZERO; digit2<=TWO; digit3<=EIGHT; end
      16'd8207: begin digit0<=SEVEN; digit1<=ZERO; digit2<=TWO; digit3<=EIGHT; end
      16'd8208: begin digit0<=EIGHT; digit1<=ZERO; digit2<=TWO; digit3<=EIGHT; end
      16'd8209: begin digit0<=NINE; digit1<=ZERO; digit2<=TWO; digit3<=EIGHT; end
      16'd8210: begin digit0<=ZERO; digit1<=ONE; digit2<=TWO; digit3<=EIGHT; end
      16'd8211: begin digit0<=ONE; digit1<=ONE; digit2<=TWO; digit3<=EIGHT; end
      16'd8212: begin digit0<=TWO; digit1<=ONE; digit2<=TWO; digit3<=EIGHT; end
      16'd8213: begin digit0<=THREE; digit1<=ONE; digit2<=TWO; digit3<=EIGHT; end
      16'd8214: begin digit0<=FOUR; digit1<=ONE; digit2<=TWO; digit3<=EIGHT; end
      16'd8215: begin digit0<=FIVE; digit1<=ONE; digit2<=TWO; digit3<=EIGHT; end
      16'd8216: begin digit0<=SIX; digit1<=ONE; digit2<=TWO; digit3<=EIGHT; end
      16'd8217: begin digit0<=SEVEN; digit1<=ONE; digit2<=TWO; digit3<=EIGHT; end
      16'd8218: begin digit0<=EIGHT; digit1<=ONE; digit2<=TWO; digit3<=EIGHT; end
      16'd8219: begin digit0<=NINE; digit1<=ONE; digit2<=TWO; digit3<=EIGHT; end
      16'd8220: begin digit0<=ZERO; digit1<=TWO; digit2<=TWO; digit3<=EIGHT; end
      16'd8221: begin digit0<=ONE; digit1<=TWO; digit2<=TWO; digit3<=EIGHT; end
      16'd8222: begin digit0<=TWO; digit1<=TWO; digit2<=TWO; digit3<=EIGHT; end
      16'd8223: begin digit0<=THREE; digit1<=TWO; digit2<=TWO; digit3<=EIGHT; end
      16'd8224: begin digit0<=FOUR; digit1<=TWO; digit2<=TWO; digit3<=EIGHT; end
      16'd8225: begin digit0<=FIVE; digit1<=TWO; digit2<=TWO; digit3<=EIGHT; end
      16'd8226: begin digit0<=SIX; digit1<=TWO; digit2<=TWO; digit3<=EIGHT; end
      16'd8227: begin digit0<=SEVEN; digit1<=TWO; digit2<=TWO; digit3<=EIGHT; end
      16'd8228: begin digit0<=EIGHT; digit1<=TWO; digit2<=TWO; digit3<=EIGHT; end
      16'd8229: begin digit0<=NINE; digit1<=TWO; digit2<=TWO; digit3<=EIGHT; end
      16'd8230: begin digit0<=ZERO; digit1<=THREE; digit2<=TWO; digit3<=EIGHT; end
      16'd8231: begin digit0<=ONE; digit1<=THREE; digit2<=TWO; digit3<=EIGHT; end
      16'd8232: begin digit0<=TWO; digit1<=THREE; digit2<=TWO; digit3<=EIGHT; end
      16'd8233: begin digit0<=THREE; digit1<=THREE; digit2<=TWO; digit3<=EIGHT; end
      16'd8234: begin digit0<=FOUR; digit1<=THREE; digit2<=TWO; digit3<=EIGHT; end
      16'd8235: begin digit0<=FIVE; digit1<=THREE; digit2<=TWO; digit3<=EIGHT; end
      16'd8236: begin digit0<=SIX; digit1<=THREE; digit2<=TWO; digit3<=EIGHT; end
      16'd8237: begin digit0<=SEVEN; digit1<=THREE; digit2<=TWO; digit3<=EIGHT; end
      16'd8238: begin digit0<=EIGHT; digit1<=THREE; digit2<=TWO; digit3<=EIGHT; end
      16'd8239: begin digit0<=NINE; digit1<=THREE; digit2<=TWO; digit3<=EIGHT; end
      16'd8240: begin digit0<=ZERO; digit1<=FOUR; digit2<=TWO; digit3<=EIGHT; end
      16'd8241: begin digit0<=ONE; digit1<=FOUR; digit2<=TWO; digit3<=EIGHT; end
      16'd8242: begin digit0<=TWO; digit1<=FOUR; digit2<=TWO; digit3<=EIGHT; end
      16'd8243: begin digit0<=THREE; digit1<=FOUR; digit2<=TWO; digit3<=EIGHT; end
      16'd8244: begin digit0<=FOUR; digit1<=FOUR; digit2<=TWO; digit3<=EIGHT; end
      16'd8245: begin digit0<=FIVE; digit1<=FOUR; digit2<=TWO; digit3<=EIGHT; end
      16'd8246: begin digit0<=SIX; digit1<=FOUR; digit2<=TWO; digit3<=EIGHT; end
      16'd8247: begin digit0<=SEVEN; digit1<=FOUR; digit2<=TWO; digit3<=EIGHT; end
      16'd8248: begin digit0<=EIGHT; digit1<=FOUR; digit2<=TWO; digit3<=EIGHT; end
      16'd8249: begin digit0<=NINE; digit1<=FOUR; digit2<=TWO; digit3<=EIGHT; end
      16'd8250: begin digit0<=ZERO; digit1<=FIVE; digit2<=TWO; digit3<=EIGHT; end
      16'd8251: begin digit0<=ONE; digit1<=FIVE; digit2<=TWO; digit3<=EIGHT; end
      16'd8252: begin digit0<=TWO; digit1<=FIVE; digit2<=TWO; digit3<=EIGHT; end
      16'd8253: begin digit0<=THREE; digit1<=FIVE; digit2<=TWO; digit3<=EIGHT; end
      16'd8254: begin digit0<=FOUR; digit1<=FIVE; digit2<=TWO; digit3<=EIGHT; end
      16'd8255: begin digit0<=FIVE; digit1<=FIVE; digit2<=TWO; digit3<=EIGHT; end
      16'd8256: begin digit0<=SIX; digit1<=FIVE; digit2<=TWO; digit3<=EIGHT; end
      16'd8257: begin digit0<=SEVEN; digit1<=FIVE; digit2<=TWO; digit3<=EIGHT; end
      16'd8258: begin digit0<=EIGHT; digit1<=FIVE; digit2<=TWO; digit3<=EIGHT; end
      16'd8259: begin digit0<=NINE; digit1<=FIVE; digit2<=TWO; digit3<=EIGHT; end
      16'd8260: begin digit0<=ZERO; digit1<=SIX; digit2<=TWO; digit3<=EIGHT; end
      16'd8261: begin digit0<=ONE; digit1<=SIX; digit2<=TWO; digit3<=EIGHT; end
      16'd8262: begin digit0<=TWO; digit1<=SIX; digit2<=TWO; digit3<=EIGHT; end
      16'd8263: begin digit0<=THREE; digit1<=SIX; digit2<=TWO; digit3<=EIGHT; end
      16'd8264: begin digit0<=FOUR; digit1<=SIX; digit2<=TWO; digit3<=EIGHT; end
      16'd8265: begin digit0<=FIVE; digit1<=SIX; digit2<=TWO; digit3<=EIGHT; end
      16'd8266: begin digit0<=SIX; digit1<=SIX; digit2<=TWO; digit3<=EIGHT; end
      16'd8267: begin digit0<=SEVEN; digit1<=SIX; digit2<=TWO; digit3<=EIGHT; end
      16'd8268: begin digit0<=EIGHT; digit1<=SIX; digit2<=TWO; digit3<=EIGHT; end
      16'd8269: begin digit0<=NINE; digit1<=SIX; digit2<=TWO; digit3<=EIGHT; end
      16'd8270: begin digit0<=ZERO; digit1<=SEVEN; digit2<=TWO; digit3<=EIGHT; end
      16'd8271: begin digit0<=ONE; digit1<=SEVEN; digit2<=TWO; digit3<=EIGHT; end
      16'd8272: begin digit0<=TWO; digit1<=SEVEN; digit2<=TWO; digit3<=EIGHT; end
      16'd8273: begin digit0<=THREE; digit1<=SEVEN; digit2<=TWO; digit3<=EIGHT; end
      16'd8274: begin digit0<=FOUR; digit1<=SEVEN; digit2<=TWO; digit3<=EIGHT; end
      16'd8275: begin digit0<=FIVE; digit1<=SEVEN; digit2<=TWO; digit3<=EIGHT; end
      16'd8276: begin digit0<=SIX; digit1<=SEVEN; digit2<=TWO; digit3<=EIGHT; end
      16'd8277: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=TWO; digit3<=EIGHT; end
      16'd8278: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=TWO; digit3<=EIGHT; end
      16'd8279: begin digit0<=NINE; digit1<=SEVEN; digit2<=TWO; digit3<=EIGHT; end
      16'd8280: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=EIGHT; end
      16'd8281: begin digit0<=ONE; digit1<=EIGHT; digit2<=TWO; digit3<=EIGHT; end
      16'd8282: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=EIGHT; end
      16'd8283: begin digit0<=THREE; digit1<=EIGHT; digit2<=TWO; digit3<=EIGHT; end
      16'd8284: begin digit0<=FOUR; digit1<=EIGHT; digit2<=TWO; digit3<=EIGHT; end
      16'd8285: begin digit0<=FIVE; digit1<=EIGHT; digit2<=TWO; digit3<=EIGHT; end
      16'd8286: begin digit0<=SIX; digit1<=EIGHT; digit2<=TWO; digit3<=EIGHT; end
      16'd8287: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=TWO; digit3<=EIGHT; end
      16'd8288: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=TWO; digit3<=EIGHT; end
      16'd8289: begin digit0<=NINE; digit1<=EIGHT; digit2<=TWO; digit3<=EIGHT; end
      16'd8290: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=EIGHT; end
      16'd8291: begin digit0<=ONE; digit1<=NINE; digit2<=TWO; digit3<=EIGHT; end
      16'd8292: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=EIGHT; end
      16'd8293: begin digit0<=THREE; digit1<=NINE; digit2<=TWO; digit3<=EIGHT; end
      16'd8294: begin digit0<=FOUR; digit1<=NINE; digit2<=TWO; digit3<=EIGHT; end
      16'd8295: begin digit0<=FIVE; digit1<=NINE; digit2<=TWO; digit3<=EIGHT; end
      16'd8296: begin digit0<=SIX; digit1<=NINE; digit2<=TWO; digit3<=EIGHT; end
      16'd8297: begin digit0<=SEVEN; digit1<=NINE; digit2<=TWO; digit3<=EIGHT; end
      16'd8298: begin digit0<=EIGHT; digit1<=NINE; digit2<=TWO; digit3<=EIGHT; end
      16'd8299: begin digit0<=NINE; digit1<=NINE; digit2<=TWO; digit3<=EIGHT; end
	  16'd8300: begin digit0<=ZERO; digit1<=ZERO; digit2<=THREE; digit3<=EIGHT; end
      16'd8301: begin digit0<=ONE; digit1<=ZERO; digit2<=THREE; digit3<=EIGHT; end
      16'd8302: begin digit0<=TWO; digit1<=ZERO; digit2<=THREE; digit3<=EIGHT; end
      16'd8303: begin digit0<=THREE; digit1<=ZERO; digit2<=THREE; digit3<=EIGHT; end
      16'd8304: begin digit0<=FOUR; digit1<=ZERO; digit2<=THREE; digit3<=EIGHT; end
      16'd8305: begin digit0<=FIVE; digit1<=ZERO; digit2<=THREE; digit3<=EIGHT; end
      16'd8306: begin digit0<=SIX; digit1<=ZERO; digit2<=THREE; digit3<=EIGHT; end
      16'd8307: begin digit0<=SEVEN; digit1<=ZERO; digit2<=THREE; digit3<=EIGHT; end
      16'd8308: begin digit0<=EIGHT; digit1<=ZERO; digit2<=THREE; digit3<=EIGHT; end
      16'd8309: begin digit0<=NINE; digit1<=ZERO; digit2<=THREE; digit3<=EIGHT; end
      16'd8310: begin digit0<=ZERO; digit1<=ONE; digit2<=THREE; digit3<=EIGHT; end
      16'd8311: begin digit0<=ONE; digit1<=ONE; digit2<=THREE; digit3<=EIGHT; end
      16'd8312: begin digit0<=TWO; digit1<=ONE; digit2<=THREE; digit3<=EIGHT; end
      16'd8313: begin digit0<=THREE; digit1<=ONE; digit2<=THREE; digit3<=EIGHT; end
      16'd8314: begin digit0<=FOUR; digit1<=ONE; digit2<=THREE; digit3<=EIGHT; end
      16'd8315: begin digit0<=FIVE; digit1<=ONE; digit2<=THREE; digit3<=EIGHT; end
      16'd8316: begin digit0<=SIX; digit1<=ONE; digit2<=THREE; digit3<=EIGHT; end
      16'd8317: begin digit0<=SEVEN; digit1<=ONE; digit2<=THREE; digit3<=EIGHT; end
      16'd8318: begin digit0<=EIGHT; digit1<=ONE; digit2<=THREE; digit3<=EIGHT; end
      16'd8319: begin digit0<=NINE; digit1<=ONE; digit2<=THREE; digit3<=EIGHT; end
      16'd8320: begin digit0<=ZERO; digit1<=TWO; digit2<=THREE; digit3<=EIGHT; end
      16'd8321: begin digit0<=ONE; digit1<=TWO; digit2<=THREE; digit3<=EIGHT; end
      16'd8322: begin digit0<=TWO; digit1<=TWO; digit2<=THREE; digit3<=EIGHT; end
      16'd8323: begin digit0<=THREE; digit1<=TWO; digit2<=THREE; digit3<=EIGHT; end
      16'd8324: begin digit0<=FOUR; digit1<=TWO; digit2<=THREE; digit3<=EIGHT; end
      16'd8325: begin digit0<=FIVE; digit1<=TWO; digit2<=THREE; digit3<=EIGHT; end
      16'd8326: begin digit0<=SIX; digit1<=TWO; digit2<=THREE; digit3<=EIGHT; end
      16'd8327: begin digit0<=SEVEN; digit1<=TWO; digit2<=THREE; digit3<=EIGHT; end
      16'd8328: begin digit0<=EIGHT; digit1<=TWO; digit2<=THREE; digit3<=EIGHT; end
      16'd8329: begin digit0<=NINE; digit1<=TWO; digit2<=THREE; digit3<=EIGHT; end
      16'd8330: begin digit0<=ZERO; digit1<=THREE; digit2<=THREE; digit3<=EIGHT; end
      16'd8331: begin digit0<=ONE; digit1<=THREE; digit2<=THREE; digit3<=EIGHT; end
      16'd8332: begin digit0<=TWO; digit1<=THREE; digit2<=THREE; digit3<=EIGHT; end
      16'd8333: begin digit0<=THREE; digit1<=THREE; digit2<=THREE; digit3<=EIGHT; end
      16'd8334: begin digit0<=FOUR; digit1<=THREE; digit2<=THREE; digit3<=EIGHT; end
      16'd8335: begin digit0<=FIVE; digit1<=THREE; digit2<=THREE; digit3<=EIGHT; end
      16'd8336: begin digit0<=SIX; digit1<=THREE; digit2<=THREE; digit3<=EIGHT; end
      16'd8337: begin digit0<=SEVEN; digit1<=THREE; digit2<=THREE; digit3<=EIGHT; end
      16'd8338: begin digit0<=EIGHT; digit1<=THREE; digit2<=THREE; digit3<=EIGHT; end
      16'd8339: begin digit0<=NINE; digit1<=THREE; digit2<=THREE; digit3<=EIGHT; end
      16'd8340: begin digit0<=ZERO; digit1<=FOUR; digit2<=THREE; digit3<=EIGHT; end
      16'd8341: begin digit0<=ONE; digit1<=FOUR; digit2<=THREE; digit3<=EIGHT; end
      16'd8342: begin digit0<=TWO; digit1<=FOUR; digit2<=THREE; digit3<=EIGHT; end
      16'd8343: begin digit0<=THREE; digit1<=FOUR; digit2<=THREE; digit3<=EIGHT; end
      16'd8344: begin digit0<=FOUR; digit1<=FOUR; digit2<=THREE; digit3<=EIGHT; end
      16'd8345: begin digit0<=FIVE; digit1<=FOUR; digit2<=THREE; digit3<=EIGHT; end
      16'd8346: begin digit0<=SIX; digit1<=FOUR; digit2<=THREE; digit3<=EIGHT; end
      16'd8347: begin digit0<=SEVEN; digit1<=FOUR; digit2<=THREE; digit3<=EIGHT; end
      16'd8348: begin digit0<=EIGHT; digit1<=FOUR; digit2<=THREE; digit3<=EIGHT; end
      16'd8349: begin digit0<=NINE; digit1<=FOUR; digit2<=THREE; digit3<=EIGHT; end
      16'd8350: begin digit0<=ZERO; digit1<=FIVE; digit2<=THREE; digit3<=EIGHT; end
      16'd8351: begin digit0<=ONE; digit1<=FIVE; digit2<=THREE; digit3<=EIGHT; end
      16'd8352: begin digit0<=TWO; digit1<=FIVE; digit2<=THREE; digit3<=EIGHT; end
      16'd8353: begin digit0<=THREE; digit1<=FIVE; digit2<=THREE; digit3<=EIGHT; end
      16'd8354: begin digit0<=FOUR; digit1<=FIVE; digit2<=THREE; digit3<=EIGHT; end
      16'd8355: begin digit0<=FIVE; digit1<=FIVE; digit2<=THREE; digit3<=EIGHT; end
      16'd8356: begin digit0<=SIX; digit1<=FIVE; digit2<=THREE; digit3<=EIGHT; end
      16'd8357: begin digit0<=SEVEN; digit1<=FIVE; digit2<=THREE; digit3<=EIGHT; end
      16'd8358: begin digit0<=EIGHT; digit1<=FIVE; digit2<=THREE; digit3<=EIGHT; end
      16'd8359: begin digit0<=NINE; digit1<=FIVE; digit2<=THREE; digit3<=EIGHT; end
      16'd8360: begin digit0<=ZERO; digit1<=SIX; digit2<=THREE; digit3<=EIGHT; end
      16'd8361: begin digit0<=ONE; digit1<=SIX; digit2<=THREE; digit3<=EIGHT; end
      16'd8362: begin digit0<=TWO; digit1<=SIX; digit2<=THREE; digit3<=EIGHT; end
      16'd8363: begin digit0<=THREE; digit1<=SIX; digit2<=THREE; digit3<=EIGHT; end
      16'd8364: begin digit0<=FOUR; digit1<=SIX; digit2<=THREE; digit3<=EIGHT; end
      16'd8365: begin digit0<=FIVE; digit1<=SIX; digit2<=THREE; digit3<=EIGHT; end
      16'd8366: begin digit0<=SIX; digit1<=SIX; digit2<=THREE; digit3<=EIGHT; end
      16'd8367: begin digit0<=SEVEN; digit1<=SIX; digit2<=THREE; digit3<=EIGHT; end
      16'd8368: begin digit0<=EIGHT; digit1<=SIX; digit2<=THREE; digit3<=EIGHT; end
      16'd8369: begin digit0<=NINE; digit1<=SIX; digit2<=THREE; digit3<=EIGHT; end
      16'd8370: begin digit0<=ZERO; digit1<=SEVEN; digit2<=THREE; digit3<=EIGHT; end
      16'd8371: begin digit0<=ONE; digit1<=SEVEN; digit2<=THREE; digit3<=EIGHT; end
      16'd8372: begin digit0<=TWO; digit1<=SEVEN; digit2<=THREE; digit3<=EIGHT; end
      16'd8373: begin digit0<=THREE; digit1<=SEVEN; digit2<=THREE; digit3<=EIGHT; end
      16'd8374: begin digit0<=FOUR; digit1<=SEVEN; digit2<=THREE; digit3<=EIGHT; end
      16'd8375: begin digit0<=FIVE; digit1<=SEVEN; digit2<=THREE; digit3<=EIGHT; end
      16'd8376: begin digit0<=SIX; digit1<=SEVEN; digit2<=THREE; digit3<=EIGHT; end
      16'd8377: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=THREE; digit3<=EIGHT; end
      16'd8378: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=THREE; digit3<=EIGHT; end
      16'd8379: begin digit0<=NINE; digit1<=SEVEN; digit2<=THREE; digit3<=EIGHT; end
      16'd8380: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=EIGHT; end
      16'd8381: begin digit0<=ONE; digit1<=EIGHT; digit2<=THREE; digit3<=EIGHT; end
      16'd8382: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=EIGHT; end
      16'd8383: begin digit0<=THREE; digit1<=EIGHT; digit2<=THREE; digit3<=EIGHT; end
      16'd8384: begin digit0<=FOUR; digit1<=EIGHT; digit2<=THREE; digit3<=EIGHT; end
      16'd8385: begin digit0<=FIVE; digit1<=EIGHT; digit2<=THREE; digit3<=EIGHT; end
      16'd8386: begin digit0<=SIX; digit1<=EIGHT; digit2<=THREE; digit3<=EIGHT; end
      16'd8387: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=THREE; digit3<=EIGHT; end
      16'd8388: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=THREE; digit3<=EIGHT; end
      16'd8389: begin digit0<=NINE; digit1<=EIGHT; digit2<=THREE; digit3<=EIGHT; end
      16'd8390: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=EIGHT; end
      16'd8391: begin digit0<=ONE; digit1<=NINE; digit2<=THREE; digit3<=EIGHT; end
      16'd8392: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=EIGHT; end
      16'd8393: begin digit0<=THREE; digit1<=NINE; digit2<=THREE; digit3<=EIGHT; end
      16'd8394: begin digit0<=FOUR; digit1<=NINE; digit2<=THREE; digit3<=EIGHT; end
      16'd8395: begin digit0<=FIVE; digit1<=NINE; digit2<=THREE; digit3<=EIGHT; end
      16'd8396: begin digit0<=SIX; digit1<=NINE; digit2<=THREE; digit3<=EIGHT; end
      16'd8397: begin digit0<=SEVEN; digit1<=NINE; digit2<=THREE; digit3<=EIGHT; end
      16'd8398: begin digit0<=EIGHT; digit1<=NINE; digit2<=THREE; digit3<=EIGHT; end
      16'd8399: begin digit0<=NINE; digit1<=NINE; digit2<=THREE; digit3<=EIGHT; end
	  16'd8400: begin digit0<=ZERO; digit1<=ZERO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8401: begin digit0<=ONE; digit1<=ZERO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8402: begin digit0<=TWO; digit1<=ZERO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8403: begin digit0<=THREE; digit1<=ZERO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8404: begin digit0<=FOUR; digit1<=ZERO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8405: begin digit0<=FIVE; digit1<=ZERO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8406: begin digit0<=SIX; digit1<=ZERO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8407: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8408: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8409: begin digit0<=NINE; digit1<=ZERO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8410: begin digit0<=ZERO; digit1<=ONE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8411: begin digit0<=ONE; digit1<=ONE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8412: begin digit0<=TWO; digit1<=ONE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8413: begin digit0<=THREE; digit1<=ONE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8414: begin digit0<=FOUR; digit1<=ONE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8415: begin digit0<=FIVE; digit1<=ONE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8416: begin digit0<=SIX; digit1<=ONE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8417: begin digit0<=SEVEN; digit1<=ONE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8418: begin digit0<=EIGHT; digit1<=ONE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8419: begin digit0<=NINE; digit1<=ONE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8420: begin digit0<=ZERO; digit1<=TWO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8421: begin digit0<=ONE; digit1<=TWO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8422: begin digit0<=TWO; digit1<=TWO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8423: begin digit0<=THREE; digit1<=TWO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8424: begin digit0<=FOUR; digit1<=TWO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8425: begin digit0<=FIVE; digit1<=TWO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8426: begin digit0<=SIX; digit1<=TWO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8427: begin digit0<=SEVEN; digit1<=TWO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8428: begin digit0<=EIGHT; digit1<=TWO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8429: begin digit0<=NINE; digit1<=TWO; digit2<=FOUR; digit3<=EIGHT; end
      16'd8430: begin digit0<=ZERO; digit1<=THREE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8431: begin digit0<=ONE; digit1<=THREE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8432: begin digit0<=TWO; digit1<=THREE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8433: begin digit0<=THREE; digit1<=THREE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8434: begin digit0<=FOUR; digit1<=THREE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8435: begin digit0<=FIVE; digit1<=THREE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8436: begin digit0<=SIX; digit1<=THREE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8437: begin digit0<=SEVEN; digit1<=THREE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8438: begin digit0<=EIGHT; digit1<=THREE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8439: begin digit0<=NINE; digit1<=THREE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8440: begin digit0<=ZERO; digit1<=FOUR; digit2<=FOUR; digit3<=EIGHT; end
      16'd8441: begin digit0<=ONE; digit1<=FOUR; digit2<=FOUR; digit3<=EIGHT; end
      16'd8442: begin digit0<=TWO; digit1<=FOUR; digit2<=FOUR; digit3<=EIGHT; end
      16'd8443: begin digit0<=THREE; digit1<=FOUR; digit2<=FOUR; digit3<=EIGHT; end
      16'd8444: begin digit0<=FOUR; digit1<=FOUR; digit2<=FOUR; digit3<=EIGHT; end
      16'd8445: begin digit0<=FIVE; digit1<=FOUR; digit2<=FOUR; digit3<=EIGHT; end
      16'd8446: begin digit0<=SIX; digit1<=FOUR; digit2<=FOUR; digit3<=EIGHT; end
      16'd8447: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FOUR; digit3<=EIGHT; end
      16'd8448: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FOUR; digit3<=EIGHT; end
      16'd8449: begin digit0<=NINE; digit1<=FOUR; digit2<=FOUR; digit3<=EIGHT; end
      16'd8450: begin digit0<=ZERO; digit1<=FIVE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8451: begin digit0<=ONE; digit1<=FIVE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8452: begin digit0<=TWO; digit1<=FIVE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8453: begin digit0<=THREE; digit1<=FIVE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8454: begin digit0<=FOUR; digit1<=FIVE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8455: begin digit0<=FIVE; digit1<=FIVE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8456: begin digit0<=SIX; digit1<=FIVE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8457: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8458: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8459: begin digit0<=NINE; digit1<=FIVE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8460: begin digit0<=ZERO; digit1<=SIX; digit2<=FOUR; digit3<=EIGHT; end
      16'd8461: begin digit0<=ONE; digit1<=SIX; digit2<=FOUR; digit3<=EIGHT; end
      16'd8462: begin digit0<=TWO; digit1<=SIX; digit2<=FOUR; digit3<=EIGHT; end
      16'd8463: begin digit0<=THREE; digit1<=SIX; digit2<=FOUR; digit3<=EIGHT; end
      16'd8464: begin digit0<=FOUR; digit1<=SIX; digit2<=FOUR; digit3<=EIGHT; end
      16'd8465: begin digit0<=FIVE; digit1<=SIX; digit2<=FOUR; digit3<=EIGHT; end
      16'd8466: begin digit0<=SIX; digit1<=SIX; digit2<=FOUR; digit3<=EIGHT; end
      16'd8467: begin digit0<=SEVEN; digit1<=SIX; digit2<=FOUR; digit3<=EIGHT; end
      16'd8468: begin digit0<=EIGHT; digit1<=SIX; digit2<=FOUR; digit3<=EIGHT; end
      16'd8469: begin digit0<=NINE; digit1<=SIX; digit2<=FOUR; digit3<=EIGHT; end
      16'd8470: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FOUR; digit3<=EIGHT; end
      16'd8471: begin digit0<=ONE; digit1<=SEVEN; digit2<=FOUR; digit3<=EIGHT; end
      16'd8472: begin digit0<=TWO; digit1<=SEVEN; digit2<=FOUR; digit3<=EIGHT; end
      16'd8473: begin digit0<=THREE; digit1<=SEVEN; digit2<=FOUR; digit3<=EIGHT; end
      16'd8474: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FOUR; digit3<=EIGHT; end
      16'd8475: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FOUR; digit3<=EIGHT; end
      16'd8476: begin digit0<=SIX; digit1<=SEVEN; digit2<=FOUR; digit3<=EIGHT; end
      16'd8477: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FOUR; digit3<=EIGHT; end
      16'd8478: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FOUR; digit3<=EIGHT; end
      16'd8479: begin digit0<=NINE; digit1<=SEVEN; digit2<=FOUR; digit3<=EIGHT; end
      16'd8480: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=EIGHT; end
      16'd8481: begin digit0<=ONE; digit1<=EIGHT; digit2<=FOUR; digit3<=EIGHT; end
      16'd8482: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=EIGHT; end
      16'd8483: begin digit0<=THREE; digit1<=EIGHT; digit2<=FOUR; digit3<=EIGHT; end
      16'd8484: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FOUR; digit3<=EIGHT; end
      16'd8485: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FOUR; digit3<=EIGHT; end
      16'd8486: begin digit0<=SIX; digit1<=EIGHT; digit2<=FOUR; digit3<=EIGHT; end
      16'd8487: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FOUR; digit3<=EIGHT; end
      16'd8488: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FOUR; digit3<=EIGHT; end
      16'd8489: begin digit0<=NINE; digit1<=EIGHT; digit2<=FOUR; digit3<=EIGHT; end
      16'd8490: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8491: begin digit0<=ONE; digit1<=NINE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8492: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8493: begin digit0<=THREE; digit1<=NINE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8494: begin digit0<=FOUR; digit1<=NINE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8495: begin digit0<=FIVE; digit1<=NINE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8496: begin digit0<=SIX; digit1<=NINE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8497: begin digit0<=SEVEN; digit1<=NINE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8498: begin digit0<=EIGHT; digit1<=NINE; digit2<=FOUR; digit3<=EIGHT; end
      16'd8499: begin digit0<=NINE; digit1<=NINE; digit2<=FOUR; digit3<=EIGHT; end
	  16'd8500: begin digit0<=ZERO; digit1<=ZERO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8501: begin digit0<=ONE; digit1<=ZERO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8502: begin digit0<=TWO; digit1<=ZERO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8503: begin digit0<=THREE; digit1<=ZERO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8504: begin digit0<=FOUR; digit1<=ZERO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8505: begin digit0<=FIVE; digit1<=ZERO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8506: begin digit0<=SIX; digit1<=ZERO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8507: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8508: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8509: begin digit0<=NINE; digit1<=ZERO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8510: begin digit0<=ZERO; digit1<=ONE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8511: begin digit0<=ONE; digit1<=ONE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8512: begin digit0<=TWO; digit1<=ONE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8513: begin digit0<=THREE; digit1<=ONE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8514: begin digit0<=FOUR; digit1<=ONE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8515: begin digit0<=FIVE; digit1<=ONE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8516: begin digit0<=SIX; digit1<=ONE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8517: begin digit0<=SEVEN; digit1<=ONE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8518: begin digit0<=EIGHT; digit1<=ONE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8519: begin digit0<=NINE; digit1<=ONE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8520: begin digit0<=ZERO; digit1<=TWO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8521: begin digit0<=ONE; digit1<=TWO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8522: begin digit0<=TWO; digit1<=TWO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8523: begin digit0<=THREE; digit1<=TWO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8524: begin digit0<=FOUR; digit1<=TWO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8525: begin digit0<=FIVE; digit1<=TWO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8526: begin digit0<=SIX; digit1<=TWO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8527: begin digit0<=SEVEN; digit1<=TWO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8528: begin digit0<=EIGHT; digit1<=TWO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8529: begin digit0<=NINE; digit1<=TWO; digit2<=FIVE; digit3<=EIGHT; end
      16'd8530: begin digit0<=ZERO; digit1<=THREE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8531: begin digit0<=ONE; digit1<=THREE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8532: begin digit0<=TWO; digit1<=THREE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8533: begin digit0<=THREE; digit1<=THREE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8534: begin digit0<=FOUR; digit1<=THREE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8535: begin digit0<=FIVE; digit1<=THREE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8536: begin digit0<=SIX; digit1<=THREE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8537: begin digit0<=SEVEN; digit1<=THREE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8538: begin digit0<=EIGHT; digit1<=THREE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8539: begin digit0<=NINE; digit1<=THREE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8540: begin digit0<=ZERO; digit1<=FOUR; digit2<=FIVE; digit3<=EIGHT; end
      16'd8541: begin digit0<=ONE; digit1<=FOUR; digit2<=FIVE; digit3<=EIGHT; end
      16'd8542: begin digit0<=TWO; digit1<=FOUR; digit2<=FIVE; digit3<=EIGHT; end
      16'd8543: begin digit0<=THREE; digit1<=FOUR; digit2<=FIVE; digit3<=EIGHT; end
      16'd8544: begin digit0<=FOUR; digit1<=FOUR; digit2<=FIVE; digit3<=EIGHT; end
      16'd8545: begin digit0<=FIVE; digit1<=FOUR; digit2<=FIVE; digit3<=EIGHT; end
      16'd8546: begin digit0<=SIX; digit1<=FOUR; digit2<=FIVE; digit3<=EIGHT; end
      16'd8547: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FIVE; digit3<=EIGHT; end
      16'd8548: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FIVE; digit3<=EIGHT; end
      16'd8549: begin digit0<=NINE; digit1<=FOUR; digit2<=FIVE; digit3<=EIGHT; end
      16'd8550: begin digit0<=ZERO; digit1<=FIVE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8551: begin digit0<=ONE; digit1<=FIVE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8552: begin digit0<=TWO; digit1<=FIVE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8553: begin digit0<=THREE; digit1<=FIVE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8554: begin digit0<=FOUR; digit1<=FIVE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8555: begin digit0<=FIVE; digit1<=FIVE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8556: begin digit0<=SIX; digit1<=FIVE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8557: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8558: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8559: begin digit0<=NINE; digit1<=FIVE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8560: begin digit0<=ZERO; digit1<=SIX; digit2<=FIVE; digit3<=EIGHT; end
      16'd8561: begin digit0<=ONE; digit1<=SIX; digit2<=FIVE; digit3<=EIGHT; end
      16'd8562: begin digit0<=TWO; digit1<=SIX; digit2<=FIVE; digit3<=EIGHT; end
      16'd8563: begin digit0<=THREE; digit1<=SIX; digit2<=FIVE; digit3<=EIGHT; end
      16'd8564: begin digit0<=FOUR; digit1<=SIX; digit2<=FIVE; digit3<=EIGHT; end
      16'd8565: begin digit0<=FIVE; digit1<=SIX; digit2<=FIVE; digit3<=EIGHT; end
      16'd8566: begin digit0<=SIX; digit1<=SIX; digit2<=FIVE; digit3<=EIGHT; end
      16'd8567: begin digit0<=SEVEN; digit1<=SIX; digit2<=FIVE; digit3<=EIGHT; end
      16'd8568: begin digit0<=EIGHT; digit1<=SIX; digit2<=FIVE; digit3<=EIGHT; end
      16'd8569: begin digit0<=NINE; digit1<=SIX; digit2<=FIVE; digit3<=EIGHT; end
      16'd8570: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FIVE; digit3<=EIGHT; end
      16'd8571: begin digit0<=ONE; digit1<=SEVEN; digit2<=FIVE; digit3<=EIGHT; end
      16'd8572: begin digit0<=TWO; digit1<=SEVEN; digit2<=FIVE; digit3<=EIGHT; end
      16'd8573: begin digit0<=THREE; digit1<=SEVEN; digit2<=FIVE; digit3<=EIGHT; end
      16'd8574: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FIVE; digit3<=EIGHT; end
      16'd8575: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FIVE; digit3<=EIGHT; end
      16'd8576: begin digit0<=SIX; digit1<=SEVEN; digit2<=FIVE; digit3<=EIGHT; end
      16'd8577: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FIVE; digit3<=EIGHT; end
      16'd8578: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FIVE; digit3<=EIGHT; end
      16'd8579: begin digit0<=NINE; digit1<=SEVEN; digit2<=FIVE; digit3<=EIGHT; end
      16'd8580: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=EIGHT; end
      16'd8581: begin digit0<=ONE; digit1<=EIGHT; digit2<=FIVE; digit3<=EIGHT; end
      16'd8582: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=EIGHT; end
      16'd8583: begin digit0<=THREE; digit1<=EIGHT; digit2<=FIVE; digit3<=EIGHT; end
      16'd8584: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FIVE; digit3<=EIGHT; end
      16'd8585: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FIVE; digit3<=EIGHT; end
      16'd8586: begin digit0<=SIX; digit1<=EIGHT; digit2<=FIVE; digit3<=EIGHT; end
      16'd8587: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FIVE; digit3<=EIGHT; end
      16'd8588: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FIVE; digit3<=EIGHT; end
      16'd8589: begin digit0<=NINE; digit1<=EIGHT; digit2<=FIVE; digit3<=EIGHT; end
      16'd8590: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8591: begin digit0<=ONE; digit1<=NINE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8592: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8593: begin digit0<=THREE; digit1<=NINE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8594: begin digit0<=FOUR; digit1<=NINE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8595: begin digit0<=FIVE; digit1<=NINE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8596: begin digit0<=SIX; digit1<=NINE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8597: begin digit0<=SEVEN; digit1<=NINE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8598: begin digit0<=EIGHT; digit1<=NINE; digit2<=FIVE; digit3<=EIGHT; end
      16'd8599: begin digit0<=NINE; digit1<=NINE; digit2<=FIVE; digit3<=EIGHT; end
	  16'd8600: begin digit0<=ZERO; digit1<=ZERO; digit2<=SIX; digit3<=EIGHT; end
      16'd8601: begin digit0<=ONE; digit1<=ZERO; digit2<=SIX; digit3<=EIGHT; end
      16'd8602: begin digit0<=TWO; digit1<=ZERO; digit2<=SIX; digit3<=EIGHT; end
      16'd8603: begin digit0<=THREE; digit1<=ZERO; digit2<=SIX; digit3<=EIGHT; end
      16'd8604: begin digit0<=FOUR; digit1<=ZERO; digit2<=SIX; digit3<=EIGHT; end
      16'd8605: begin digit0<=FIVE; digit1<=ZERO; digit2<=SIX; digit3<=EIGHT; end
      16'd8606: begin digit0<=SIX; digit1<=ZERO; digit2<=SIX; digit3<=EIGHT; end
      16'd8607: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SIX; digit3<=EIGHT; end
      16'd8608: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SIX; digit3<=EIGHT; end
      16'd8609: begin digit0<=NINE; digit1<=ZERO; digit2<=SIX; digit3<=EIGHT; end
      16'd8610: begin digit0<=ZERO; digit1<=ONE; digit2<=SIX; digit3<=EIGHT; end
      16'd8611: begin digit0<=ONE; digit1<=ONE; digit2<=SIX; digit3<=EIGHT; end
      16'd8612: begin digit0<=TWO; digit1<=ONE; digit2<=SIX; digit3<=EIGHT; end
      16'd8613: begin digit0<=THREE; digit1<=ONE; digit2<=SIX; digit3<=EIGHT; end
      16'd8614: begin digit0<=FOUR; digit1<=ONE; digit2<=SIX; digit3<=EIGHT; end
      16'd8615: begin digit0<=FIVE; digit1<=ONE; digit2<=SIX; digit3<=EIGHT; end
      16'd8616: begin digit0<=SIX; digit1<=ONE; digit2<=SIX; digit3<=EIGHT; end
      16'd8617: begin digit0<=SEVEN; digit1<=ONE; digit2<=SIX; digit3<=EIGHT; end
      16'd8618: begin digit0<=EIGHT; digit1<=ONE; digit2<=SIX; digit3<=EIGHT; end
      16'd8619: begin digit0<=NINE; digit1<=ONE; digit2<=SIX; digit3<=EIGHT; end
      16'd8620: begin digit0<=ZERO; digit1<=TWO; digit2<=SIX; digit3<=EIGHT; end
      16'd8621: begin digit0<=ONE; digit1<=TWO; digit2<=SIX; digit3<=EIGHT; end
      16'd8622: begin digit0<=TWO; digit1<=TWO; digit2<=SIX; digit3<=EIGHT; end
      16'd8623: begin digit0<=THREE; digit1<=TWO; digit2<=SIX; digit3<=EIGHT; end
      16'd8624: begin digit0<=FOUR; digit1<=TWO; digit2<=SIX; digit3<=EIGHT; end
      16'd8625: begin digit0<=FIVE; digit1<=TWO; digit2<=SIX; digit3<=EIGHT; end
      16'd8626: begin digit0<=SIX; digit1<=TWO; digit2<=SIX; digit3<=EIGHT; end
      16'd8627: begin digit0<=SEVEN; digit1<=TWO; digit2<=SIX; digit3<=EIGHT; end
      16'd8628: begin digit0<=EIGHT; digit1<=TWO; digit2<=SIX; digit3<=EIGHT; end
      16'd8629: begin digit0<=NINE; digit1<=TWO; digit2<=SIX; digit3<=EIGHT; end
      16'd8630: begin digit0<=ZERO; digit1<=THREE; digit2<=SIX; digit3<=EIGHT; end
      16'd8631: begin digit0<=ONE; digit1<=THREE; digit2<=SIX; digit3<=EIGHT; end
      16'd8632: begin digit0<=TWO; digit1<=THREE; digit2<=SIX; digit3<=EIGHT; end
      16'd8633: begin digit0<=THREE; digit1<=THREE; digit2<=SIX; digit3<=EIGHT; end
      16'd8634: begin digit0<=FOUR; digit1<=THREE; digit2<=SIX; digit3<=EIGHT; end
      16'd8635: begin digit0<=FIVE; digit1<=THREE; digit2<=SIX; digit3<=EIGHT; end
      16'd8636: begin digit0<=SIX; digit1<=THREE; digit2<=SIX; digit3<=EIGHT; end
      16'd8637: begin digit0<=SEVEN; digit1<=THREE; digit2<=SIX; digit3<=EIGHT; end
      16'd8638: begin digit0<=EIGHT; digit1<=THREE; digit2<=SIX; digit3<=EIGHT; end
      16'd8639: begin digit0<=NINE; digit1<=THREE; digit2<=SIX; digit3<=EIGHT; end
      16'd8640: begin digit0<=ZERO; digit1<=FOUR; digit2<=SIX; digit3<=EIGHT; end
      16'd8641: begin digit0<=ONE; digit1<=FOUR; digit2<=SIX; digit3<=EIGHT; end
      16'd8642: begin digit0<=TWO; digit1<=FOUR; digit2<=SIX; digit3<=EIGHT; end
      16'd8643: begin digit0<=THREE; digit1<=FOUR; digit2<=SIX; digit3<=EIGHT; end
      16'd8644: begin digit0<=FOUR; digit1<=FOUR; digit2<=SIX; digit3<=EIGHT; end
      16'd8645: begin digit0<=FIVE; digit1<=FOUR; digit2<=SIX; digit3<=EIGHT; end
      16'd8646: begin digit0<=SIX; digit1<=FOUR; digit2<=SIX; digit3<=EIGHT; end
      16'd8647: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SIX; digit3<=EIGHT; end
      16'd8648: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SIX; digit3<=EIGHT; end
      16'd8649: begin digit0<=NINE; digit1<=FOUR; digit2<=SIX; digit3<=EIGHT; end
      16'd8650: begin digit0<=ZERO; digit1<=FIVE; digit2<=SIX; digit3<=EIGHT; end
      16'd8651: begin digit0<=ONE; digit1<=FIVE; digit2<=SIX; digit3<=EIGHT; end
      16'd8652: begin digit0<=TWO; digit1<=FIVE; digit2<=SIX; digit3<=EIGHT; end
      16'd8653: begin digit0<=THREE; digit1<=FIVE; digit2<=SIX; digit3<=EIGHT; end
      16'd8654: begin digit0<=FOUR; digit1<=FIVE; digit2<=SIX; digit3<=EIGHT; end
      16'd8655: begin digit0<=FIVE; digit1<=FIVE; digit2<=SIX; digit3<=EIGHT; end
      16'd8656: begin digit0<=SIX; digit1<=FIVE; digit2<=SIX; digit3<=EIGHT; end
      16'd8657: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SIX; digit3<=EIGHT; end
      16'd8658: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SIX; digit3<=EIGHT; end
      16'd8659: begin digit0<=NINE; digit1<=FIVE; digit2<=SIX; digit3<=EIGHT; end
      16'd8660: begin digit0<=ZERO; digit1<=SIX; digit2<=SIX; digit3<=EIGHT; end
      16'd8661: begin digit0<=ONE; digit1<=SIX; digit2<=SIX; digit3<=EIGHT; end
      16'd8662: begin digit0<=TWO; digit1<=SIX; digit2<=SIX; digit3<=EIGHT; end
      16'd8663: begin digit0<=THREE; digit1<=SIX; digit2<=SIX; digit3<=EIGHT; end
      16'd8664: begin digit0<=FOUR; digit1<=SIX; digit2<=SIX; digit3<=EIGHT; end
      16'd8665: begin digit0<=FIVE; digit1<=SIX; digit2<=SIX; digit3<=EIGHT; end
      16'd8666: begin digit0<=SIX; digit1<=SIX; digit2<=SIX; digit3<=EIGHT; end
      16'd8667: begin digit0<=SEVEN; digit1<=SIX; digit2<=SIX; digit3<=EIGHT; end
      16'd8668: begin digit0<=EIGHT; digit1<=SIX; digit2<=SIX; digit3<=EIGHT; end
      16'd8669: begin digit0<=NINE; digit1<=SIX; digit2<=SIX; digit3<=EIGHT; end
      16'd8670: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SIX; digit3<=EIGHT; end
      16'd8671: begin digit0<=ONE; digit1<=SEVEN; digit2<=SIX; digit3<=EIGHT; end
      16'd8672: begin digit0<=TWO; digit1<=SEVEN; digit2<=SIX; digit3<=EIGHT; end
      16'd8673: begin digit0<=THREE; digit1<=SEVEN; digit2<=SIX; digit3<=EIGHT; end
      16'd8674: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SIX; digit3<=EIGHT; end
      16'd8675: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SIX; digit3<=EIGHT; end
      16'd8676: begin digit0<=SIX; digit1<=SEVEN; digit2<=SIX; digit3<=EIGHT; end
      16'd8677: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SIX; digit3<=EIGHT; end
      16'd8678: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SIX; digit3<=EIGHT; end
      16'd8679: begin digit0<=NINE; digit1<=SEVEN; digit2<=SIX; digit3<=EIGHT; end
      16'd8680: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=EIGHT; end
      16'd8681: begin digit0<=ONE; digit1<=EIGHT; digit2<=SIX; digit3<=EIGHT; end
      16'd8682: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=EIGHT; end
      16'd8683: begin digit0<=THREE; digit1<=EIGHT; digit2<=SIX; digit3<=EIGHT; end
      16'd8684: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SIX; digit3<=EIGHT; end
      16'd8685: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SIX; digit3<=EIGHT; end
      16'd8686: begin digit0<=SIX; digit1<=EIGHT; digit2<=SIX; digit3<=EIGHT; end
      16'd8687: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SIX; digit3<=EIGHT; end
      16'd8688: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SIX; digit3<=EIGHT; end
      16'd8689: begin digit0<=NINE; digit1<=EIGHT; digit2<=SIX; digit3<=EIGHT; end
      16'd8690: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=EIGHT; end
      16'd8691: begin digit0<=ONE; digit1<=NINE; digit2<=SIX; digit3<=EIGHT; end
      16'd8692: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=EIGHT; end
      16'd8693: begin digit0<=THREE; digit1<=NINE; digit2<=SIX; digit3<=EIGHT; end
      16'd8694: begin digit0<=FOUR; digit1<=NINE; digit2<=SIX; digit3<=EIGHT; end
      16'd8695: begin digit0<=FIVE; digit1<=NINE; digit2<=SIX; digit3<=EIGHT; end
      16'd8696: begin digit0<=SIX; digit1<=NINE; digit2<=SIX; digit3<=EIGHT; end
      16'd8697: begin digit0<=SEVEN; digit1<=NINE; digit2<=SIX; digit3<=EIGHT; end
      16'd8698: begin digit0<=EIGHT; digit1<=NINE; digit2<=SIX; digit3<=EIGHT; end
      16'd8699: begin digit0<=NINE; digit1<=NINE; digit2<=SIX; digit3<=EIGHT; end
	  16'd8700: begin digit0<=ZERO; digit1<=ZERO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8701: begin digit0<=ONE; digit1<=ZERO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8702: begin digit0<=TWO; digit1<=ZERO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8703: begin digit0<=THREE; digit1<=ZERO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8704: begin digit0<=FOUR; digit1<=ZERO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8705: begin digit0<=FIVE; digit1<=ZERO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8706: begin digit0<=SIX; digit1<=ZERO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8707: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8708: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8709: begin digit0<=NINE; digit1<=ZERO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8710: begin digit0<=ZERO; digit1<=ONE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8711: begin digit0<=ONE; digit1<=ONE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8712: begin digit0<=TWO; digit1<=ONE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8713: begin digit0<=THREE; digit1<=ONE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8714: begin digit0<=FOUR; digit1<=ONE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8715: begin digit0<=FIVE; digit1<=ONE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8716: begin digit0<=SIX; digit1<=ONE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8717: begin digit0<=SEVEN; digit1<=ONE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8718: begin digit0<=EIGHT; digit1<=ONE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8719: begin digit0<=NINE; digit1<=ONE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8720: begin digit0<=ZERO; digit1<=TWO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8721: begin digit0<=ONE; digit1<=TWO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8722: begin digit0<=TWO; digit1<=TWO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8723: begin digit0<=THREE; digit1<=TWO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8724: begin digit0<=FOUR; digit1<=TWO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8725: begin digit0<=FIVE; digit1<=TWO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8726: begin digit0<=SIX; digit1<=TWO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8727: begin digit0<=SEVEN; digit1<=TWO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8728: begin digit0<=EIGHT; digit1<=TWO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8729: begin digit0<=NINE; digit1<=TWO; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8730: begin digit0<=ZERO; digit1<=THREE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8731: begin digit0<=ONE; digit1<=THREE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8732: begin digit0<=TWO; digit1<=THREE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8733: begin digit0<=THREE; digit1<=THREE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8734: begin digit0<=FOUR; digit1<=THREE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8735: begin digit0<=FIVE; digit1<=THREE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8736: begin digit0<=SIX; digit1<=THREE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8737: begin digit0<=SEVEN; digit1<=THREE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8738: begin digit0<=EIGHT; digit1<=THREE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8739: begin digit0<=NINE; digit1<=THREE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8740: begin digit0<=ZERO; digit1<=FOUR; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8741: begin digit0<=ONE; digit1<=FOUR; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8742: begin digit0<=TWO; digit1<=FOUR; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8743: begin digit0<=THREE; digit1<=FOUR; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8744: begin digit0<=FOUR; digit1<=FOUR; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8745: begin digit0<=FIVE; digit1<=FOUR; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8746: begin digit0<=SIX; digit1<=FOUR; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8747: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8748: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8749: begin digit0<=NINE; digit1<=FOUR; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8750: begin digit0<=ZERO; digit1<=FIVE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8751: begin digit0<=ONE; digit1<=FIVE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8752: begin digit0<=TWO; digit1<=FIVE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8753: begin digit0<=THREE; digit1<=FIVE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8754: begin digit0<=FOUR; digit1<=FIVE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8755: begin digit0<=FIVE; digit1<=FIVE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8756: begin digit0<=SIX; digit1<=FIVE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8757: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8758: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8759: begin digit0<=NINE; digit1<=FIVE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8760: begin digit0<=ZERO; digit1<=SIX; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8761: begin digit0<=ONE; digit1<=SIX; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8762: begin digit0<=TWO; digit1<=SIX; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8763: begin digit0<=THREE; digit1<=SIX; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8764: begin digit0<=FOUR; digit1<=SIX; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8765: begin digit0<=FIVE; digit1<=SIX; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8766: begin digit0<=SIX; digit1<=SIX; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8767: begin digit0<=SEVEN; digit1<=SIX; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8768: begin digit0<=EIGHT; digit1<=SIX; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8769: begin digit0<=NINE; digit1<=SIX; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8770: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8771: begin digit0<=ONE; digit1<=SEVEN; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8772: begin digit0<=TWO; digit1<=SEVEN; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8773: begin digit0<=THREE; digit1<=SEVEN; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8774: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8775: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8776: begin digit0<=SIX; digit1<=SEVEN; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8777: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8778: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8779: begin digit0<=NINE; digit1<=SEVEN; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8780: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8781: begin digit0<=ONE; digit1<=EIGHT; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8782: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8783: begin digit0<=THREE; digit1<=EIGHT; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8784: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8785: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8786: begin digit0<=SIX; digit1<=EIGHT; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8787: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8788: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8789: begin digit0<=NINE; digit1<=EIGHT; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8790: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8791: begin digit0<=ONE; digit1<=NINE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8792: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8793: begin digit0<=THREE; digit1<=NINE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8794: begin digit0<=FOUR; digit1<=NINE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8795: begin digit0<=FIVE; digit1<=NINE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8796: begin digit0<=SIX; digit1<=NINE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8797: begin digit0<=SEVEN; digit1<=NINE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8798: begin digit0<=EIGHT; digit1<=NINE; digit2<=SEVEN; digit3<=EIGHT; end
      16'd8799: begin digit0<=NINE; digit1<=NINE; digit2<=SEVEN; digit3<=EIGHT; end
	  16'd8800: begin digit0<=ZERO; digit1<=ZERO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8801: begin digit0<=ONE; digit1<=ZERO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8802: begin digit0<=TWO; digit1<=ZERO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8803: begin digit0<=THREE; digit1<=ZERO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8804: begin digit0<=FOUR; digit1<=ZERO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8805: begin digit0<=FIVE; digit1<=ZERO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8806: begin digit0<=SIX; digit1<=ZERO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8807: begin digit0<=SEVEN; digit1<=ZERO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8808: begin digit0<=EIGHT; digit1<=ZERO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8809: begin digit0<=NINE; digit1<=ZERO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8810: begin digit0<=ZERO; digit1<=ONE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8811: begin digit0<=ONE; digit1<=ONE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8812: begin digit0<=TWO; digit1<=ONE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8813: begin digit0<=THREE; digit1<=ONE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8814: begin digit0<=FOUR; digit1<=ONE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8815: begin digit0<=FIVE; digit1<=ONE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8816: begin digit0<=SIX; digit1<=ONE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8817: begin digit0<=SEVEN; digit1<=ONE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8818: begin digit0<=EIGHT; digit1<=ONE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8819: begin digit0<=NINE; digit1<=ONE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8820: begin digit0<=ZERO; digit1<=TWO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8821: begin digit0<=ONE; digit1<=TWO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8822: begin digit0<=TWO; digit1<=TWO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8823: begin digit0<=THREE; digit1<=TWO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8824: begin digit0<=FOUR; digit1<=TWO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8825: begin digit0<=FIVE; digit1<=TWO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8826: begin digit0<=SIX; digit1<=TWO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8827: begin digit0<=SEVEN; digit1<=TWO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8828: begin digit0<=EIGHT; digit1<=TWO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8829: begin digit0<=NINE; digit1<=TWO; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8830: begin digit0<=ZERO; digit1<=THREE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8831: begin digit0<=ONE; digit1<=THREE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8832: begin digit0<=TWO; digit1<=THREE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8833: begin digit0<=THREE; digit1<=THREE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8834: begin digit0<=FOUR; digit1<=THREE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8835: begin digit0<=FIVE; digit1<=THREE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8836: begin digit0<=SIX; digit1<=THREE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8837: begin digit0<=SEVEN; digit1<=THREE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8838: begin digit0<=EIGHT; digit1<=THREE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8839: begin digit0<=NINE; digit1<=THREE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8840: begin digit0<=ZERO; digit1<=FOUR; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8841: begin digit0<=ONE; digit1<=FOUR; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8842: begin digit0<=TWO; digit1<=FOUR; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8843: begin digit0<=THREE; digit1<=FOUR; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8844: begin digit0<=FOUR; digit1<=FOUR; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8845: begin digit0<=FIVE; digit1<=FOUR; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8846: begin digit0<=SIX; digit1<=FOUR; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8847: begin digit0<=SEVEN; digit1<=FOUR; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8848: begin digit0<=EIGHT; digit1<=FOUR; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8849: begin digit0<=NINE; digit1<=FOUR; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8850: begin digit0<=ZERO; digit1<=FIVE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8851: begin digit0<=ONE; digit1<=FIVE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8852: begin digit0<=TWO; digit1<=FIVE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8853: begin digit0<=THREE; digit1<=FIVE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8854: begin digit0<=FOUR; digit1<=FIVE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8855: begin digit0<=FIVE; digit1<=FIVE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8856: begin digit0<=SIX; digit1<=FIVE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8857: begin digit0<=SEVEN; digit1<=FIVE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8858: begin digit0<=EIGHT; digit1<=FIVE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8859: begin digit0<=NINE; digit1<=FIVE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8860: begin digit0<=ZERO; digit1<=SIX; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8861: begin digit0<=ONE; digit1<=SIX; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8862: begin digit0<=TWO; digit1<=SIX; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8863: begin digit0<=THREE; digit1<=SIX; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8864: begin digit0<=FOUR; digit1<=SIX; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8865: begin digit0<=FIVE; digit1<=SIX; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8866: begin digit0<=SIX; digit1<=SIX; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8867: begin digit0<=SEVEN; digit1<=SIX; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8868: begin digit0<=EIGHT; digit1<=SIX; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8869: begin digit0<=NINE; digit1<=SIX; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8870: begin digit0<=ZERO; digit1<=SEVEN; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8871: begin digit0<=ONE; digit1<=SEVEN; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8872: begin digit0<=TWO; digit1<=SEVEN; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8873: begin digit0<=THREE; digit1<=SEVEN; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8874: begin digit0<=FOUR; digit1<=SEVEN; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8875: begin digit0<=FIVE; digit1<=SEVEN; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8876: begin digit0<=SIX; digit1<=SEVEN; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8877: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8878: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8879: begin digit0<=NINE; digit1<=SEVEN; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8880: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8881: begin digit0<=ONE; digit1<=EIGHT; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8882: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8883: begin digit0<=THREE; digit1<=EIGHT; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8884: begin digit0<=FOUR; digit1<=EIGHT; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8885: begin digit0<=FIVE; digit1<=EIGHT; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8886: begin digit0<=SIX; digit1<=EIGHT; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8887: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8888: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8889: begin digit0<=NINE; digit1<=EIGHT; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8890: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8891: begin digit0<=ONE; digit1<=NINE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8892: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8893: begin digit0<=THREE; digit1<=NINE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8894: begin digit0<=FOUR; digit1<=NINE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8895: begin digit0<=FIVE; digit1<=NINE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8896: begin digit0<=SIX; digit1<=NINE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8897: begin digit0<=SEVEN; digit1<=NINE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8898: begin digit0<=EIGHT; digit1<=NINE; digit2<=EIGHT; digit3<=EIGHT; end
      16'd8899: begin digit0<=NINE; digit1<=NINE; digit2<=EIGHT; digit3<=EIGHT; end
	  16'd8900: begin digit0<=ZERO; digit1<=ZERO; digit2<=NINE; digit3<=EIGHT; end
      16'd8901: begin digit0<=ONE; digit1<=ZERO; digit2<=NINE; digit3<=EIGHT; end
      16'd8902: begin digit0<=TWO; digit1<=ZERO; digit2<=NINE; digit3<=EIGHT; end
      16'd8903: begin digit0<=THREE; digit1<=ZERO; digit2<=NINE; digit3<=EIGHT; end
      16'd8904: begin digit0<=FOUR; digit1<=ZERO; digit2<=NINE; digit3<=EIGHT; end
      16'd8905: begin digit0<=FIVE; digit1<=ZERO; digit2<=NINE; digit3<=EIGHT; end
      16'd8906: begin digit0<=SIX; digit1<=ZERO; digit2<=NINE; digit3<=EIGHT; end
      16'd8907: begin digit0<=SEVEN; digit1<=ZERO; digit2<=NINE; digit3<=EIGHT; end
      16'd8908: begin digit0<=EIGHT; digit1<=ZERO; digit2<=NINE; digit3<=EIGHT; end
      16'd8909: begin digit0<=NINE; digit1<=ZERO; digit2<=NINE; digit3<=EIGHT; end
      16'd8910: begin digit0<=ZERO; digit1<=ONE; digit2<=NINE; digit3<=EIGHT; end
      16'd8911: begin digit0<=ONE; digit1<=ONE; digit2<=NINE; digit3<=EIGHT; end
      16'd8912: begin digit0<=TWO; digit1<=ONE; digit2<=NINE; digit3<=EIGHT; end
      16'd8913: begin digit0<=THREE; digit1<=ONE; digit2<=NINE; digit3<=EIGHT; end
      16'd8914: begin digit0<=FOUR; digit1<=ONE; digit2<=NINE; digit3<=EIGHT; end
      16'd8915: begin digit0<=FIVE; digit1<=ONE; digit2<=NINE; digit3<=EIGHT; end
      16'd8916: begin digit0<=SIX; digit1<=ONE; digit2<=NINE; digit3<=EIGHT; end
      16'd8917: begin digit0<=SEVEN; digit1<=ONE; digit2<=NINE; digit3<=EIGHT; end
      16'd8918: begin digit0<=EIGHT; digit1<=ONE; digit2<=NINE; digit3<=EIGHT; end
      16'd8919: begin digit0<=NINE; digit1<=ONE; digit2<=NINE; digit3<=EIGHT; end
      16'd8920: begin digit0<=ZERO; digit1<=TWO; digit2<=NINE; digit3<=EIGHT; end
      16'd8921: begin digit0<=ONE; digit1<=TWO; digit2<=NINE; digit3<=EIGHT; end
      16'd8922: begin digit0<=TWO; digit1<=TWO; digit2<=NINE; digit3<=EIGHT; end
      16'd8923: begin digit0<=THREE; digit1<=TWO; digit2<=NINE; digit3<=EIGHT; end
      16'd8924: begin digit0<=FOUR; digit1<=TWO; digit2<=NINE; digit3<=EIGHT; end
      16'd8925: begin digit0<=FIVE; digit1<=TWO; digit2<=NINE; digit3<=EIGHT; end
      16'd8926: begin digit0<=SIX; digit1<=TWO; digit2<=NINE; digit3<=EIGHT; end
      16'd8927: begin digit0<=SEVEN; digit1<=TWO; digit2<=NINE; digit3<=EIGHT; end
      16'd8928: begin digit0<=EIGHT; digit1<=TWO; digit2<=NINE; digit3<=EIGHT; end
      16'd8929: begin digit0<=NINE; digit1<=TWO; digit2<=NINE; digit3<=EIGHT; end
      16'd8930: begin digit0<=ZERO; digit1<=THREE; digit2<=NINE; digit3<=EIGHT; end
      16'd8931: begin digit0<=ONE; digit1<=THREE; digit2<=NINE; digit3<=EIGHT; end
      16'd8932: begin digit0<=TWO; digit1<=THREE; digit2<=NINE; digit3<=EIGHT; end
      16'd8933: begin digit0<=THREE; digit1<=THREE; digit2<=NINE; digit3<=EIGHT; end
      16'd8934: begin digit0<=FOUR; digit1<=THREE; digit2<=NINE; digit3<=EIGHT; end
      16'd8935: begin digit0<=FIVE; digit1<=THREE; digit2<=NINE; digit3<=EIGHT; end
      16'd8936: begin digit0<=SIX; digit1<=THREE; digit2<=NINE; digit3<=EIGHT; end
      16'd8937: begin digit0<=SEVEN; digit1<=THREE; digit2<=NINE; digit3<=EIGHT; end
      16'd8938: begin digit0<=EIGHT; digit1<=THREE; digit2<=NINE; digit3<=EIGHT; end
      16'd8939: begin digit0<=NINE; digit1<=THREE; digit2<=NINE; digit3<=EIGHT; end
      16'd8940: begin digit0<=ZERO; digit1<=FOUR; digit2<=NINE; digit3<=EIGHT; end
      16'd8941: begin digit0<=ONE; digit1<=FOUR; digit2<=NINE; digit3<=EIGHT; end
      16'd8942: begin digit0<=TWO; digit1<=FOUR; digit2<=NINE; digit3<=EIGHT; end
      16'd8943: begin digit0<=THREE; digit1<=FOUR; digit2<=NINE; digit3<=EIGHT; end
      16'd8944: begin digit0<=FOUR; digit1<=FOUR; digit2<=NINE; digit3<=EIGHT; end
      16'd8945: begin digit0<=FIVE; digit1<=FOUR; digit2<=NINE; digit3<=EIGHT; end
      16'd8946: begin digit0<=SIX; digit1<=FOUR; digit2<=NINE; digit3<=EIGHT; end
      16'd8947: begin digit0<=SEVEN; digit1<=FOUR; digit2<=NINE; digit3<=EIGHT; end
      16'd8948: begin digit0<=EIGHT; digit1<=FOUR; digit2<=NINE; digit3<=EIGHT; end
      16'd8949: begin digit0<=NINE; digit1<=FOUR; digit2<=NINE; digit3<=EIGHT; end
      16'd8950: begin digit0<=ZERO; digit1<=FIVE; digit2<=NINE; digit3<=EIGHT; end
      16'd8951: begin digit0<=ONE; digit1<=FIVE; digit2<=NINE; digit3<=EIGHT; end
      16'd8952: begin digit0<=TWO; digit1<=FIVE; digit2<=NINE; digit3<=EIGHT; end
      16'd8953: begin digit0<=THREE; digit1<=FIVE; digit2<=NINE; digit3<=EIGHT; end
      16'd8954: begin digit0<=FOUR; digit1<=FIVE; digit2<=NINE; digit3<=EIGHT; end
      16'd8955: begin digit0<=FIVE; digit1<=FIVE; digit2<=NINE; digit3<=EIGHT; end
      16'd8956: begin digit0<=SIX; digit1<=FIVE; digit2<=NINE; digit3<=EIGHT; end
      16'd8957: begin digit0<=SEVEN; digit1<=FIVE; digit2<=NINE; digit3<=EIGHT; end
      16'd8958: begin digit0<=EIGHT; digit1<=FIVE; digit2<=NINE; digit3<=EIGHT; end
      16'd8959: begin digit0<=NINE; digit1<=FIVE; digit2<=NINE; digit3<=EIGHT; end
      16'd8960: begin digit0<=ZERO; digit1<=SIX; digit2<=NINE; digit3<=EIGHT; end
      16'd8961: begin digit0<=ONE; digit1<=SIX; digit2<=NINE; digit3<=EIGHT; end
      16'd8962: begin digit0<=TWO; digit1<=SIX; digit2<=NINE; digit3<=EIGHT; end
      16'd8963: begin digit0<=THREE; digit1<=SIX; digit2<=NINE; digit3<=EIGHT; end
      16'd8964: begin digit0<=FOUR; digit1<=SIX; digit2<=NINE; digit3<=EIGHT; end
      16'd8965: begin digit0<=FIVE; digit1<=SIX; digit2<=NINE; digit3<=EIGHT; end
      16'd8966: begin digit0<=SIX; digit1<=SIX; digit2<=NINE; digit3<=EIGHT; end
      16'd8967: begin digit0<=SEVEN; digit1<=SIX; digit2<=NINE; digit3<=EIGHT; end
      16'd8968: begin digit0<=EIGHT; digit1<=SIX; digit2<=NINE; digit3<=EIGHT; end
      16'd8969: begin digit0<=NINE; digit1<=SIX; digit2<=NINE; digit3<=EIGHT; end
      16'd8970: begin digit0<=ZERO; digit1<=SEVEN; digit2<=NINE; digit3<=EIGHT; end
      16'd8971: begin digit0<=ONE; digit1<=SEVEN; digit2<=NINE; digit3<=EIGHT; end
      16'd8972: begin digit0<=TWO; digit1<=SEVEN; digit2<=NINE; digit3<=EIGHT; end
      16'd8973: begin digit0<=THREE; digit1<=SEVEN; digit2<=NINE; digit3<=EIGHT; end
      16'd8974: begin digit0<=FOUR; digit1<=SEVEN; digit2<=NINE; digit3<=EIGHT; end
      16'd8975: begin digit0<=FIVE; digit1<=SEVEN; digit2<=NINE; digit3<=EIGHT; end
      16'd8976: begin digit0<=SIX; digit1<=SEVEN; digit2<=NINE; digit3<=EIGHT; end
      16'd8977: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=NINE; digit3<=EIGHT; end
      16'd8978: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=NINE; digit3<=EIGHT; end
      16'd8979: begin digit0<=NINE; digit1<=SEVEN; digit2<=NINE; digit3<=EIGHT; end
      16'd8980: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=EIGHT; end
      16'd8981: begin digit0<=ONE; digit1<=EIGHT; digit2<=NINE; digit3<=EIGHT; end
      16'd8982: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=EIGHT; end
      16'd8983: begin digit0<=THREE; digit1<=EIGHT; digit2<=NINE; digit3<=EIGHT; end
      16'd8984: begin digit0<=FOUR; digit1<=EIGHT; digit2<=NINE; digit3<=EIGHT; end
      16'd8985: begin digit0<=FIVE; digit1<=EIGHT; digit2<=NINE; digit3<=EIGHT; end
      16'd8986: begin digit0<=SIX; digit1<=EIGHT; digit2<=NINE; digit3<=EIGHT; end
      16'd8987: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=NINE; digit3<=EIGHT; end
      16'd8988: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=NINE; digit3<=EIGHT; end
      16'd8989: begin digit0<=NINE; digit1<=EIGHT; digit2<=NINE; digit3<=EIGHT; end
      16'd8990: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=EIGHT; end
      16'd8991: begin digit0<=ONE; digit1<=NINE; digit2<=NINE; digit3<=EIGHT; end
      16'd8992: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=EIGHT; end
      16'd8993: begin digit0<=THREE; digit1<=NINE; digit2<=NINE; digit3<=EIGHT; end
      16'd8994: begin digit0<=FOUR; digit1<=NINE; digit2<=NINE; digit3<=EIGHT; end
      16'd8995: begin digit0<=FIVE; digit1<=NINE; digit2<=NINE; digit3<=EIGHT; end
      16'd8996: begin digit0<=SIX; digit1<=NINE; digit2<=NINE; digit3<=EIGHT; end
      16'd8997: begin digit0<=SEVEN; digit1<=NINE; digit2<=NINE; digit3<=EIGHT; end
      16'd8998: begin digit0<=EIGHT; digit1<=NINE; digit2<=NINE; digit3<=EIGHT; end
      16'd8999: begin digit0<=NINE; digit1<=NINE; digit2<=NINE; digit3<=EIGHT; end
	  16'd9000: begin digit0<=ZERO; digit1<=ZERO; digit2<=ZERO; digit3<=NINE; end
      16'd9001: begin digit0<=ONE; digit1<=ZERO; digit2<=ZERO; digit3<=NINE; end
      16'd9002: begin digit0<=TWO; digit1<=ZERO; digit2<=ZERO; digit3<=NINE; end
      16'd9003: begin digit0<=THREE; digit1<=ZERO; digit2<=ZERO; digit3<=NINE; end
      16'd9004: begin digit0<=FOUR; digit1<=ZERO; digit2<=ZERO; digit3<=NINE; end
      16'd9005: begin digit0<=FIVE; digit1<=ZERO; digit2<=ZERO; digit3<=NINE; end
      16'd9006: begin digit0<=SIX; digit1<=ZERO; digit2<=ZERO; digit3<=NINE; end
      16'd9007: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ZERO; digit3<=NINE; end
      16'd9008: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ZERO; digit3<=NINE; end
      16'd9009: begin digit0<=NINE; digit1<=ZERO; digit2<=ZERO; digit3<=NINE; end
      16'd9010: begin digit0<=ZERO; digit1<=ONE; digit2<=ZERO; digit3<=NINE; end
      16'd9011: begin digit0<=ONE; digit1<=ONE; digit2<=ZERO; digit3<=NINE; end
      16'd9012: begin digit0<=TWO; digit1<=ONE; digit2<=ZERO; digit3<=NINE; end
      16'd9013: begin digit0<=THREE; digit1<=ONE; digit2<=ZERO; digit3<=NINE; end
      16'd9014: begin digit0<=FOUR; digit1<=ONE; digit2<=ZERO; digit3<=NINE; end
      16'd9015: begin digit0<=FIVE; digit1<=ONE; digit2<=ZERO; digit3<=NINE; end
      16'd9016: begin digit0<=SIX; digit1<=ONE; digit2<=ZERO; digit3<=NINE; end
      16'd9017: begin digit0<=SEVEN; digit1<=ONE; digit2<=ZERO; digit3<=NINE; end
      16'd9018: begin digit0<=EIGHT; digit1<=ONE; digit2<=ZERO; digit3<=NINE; end
      16'd9019: begin digit0<=NINE; digit1<=ONE; digit2<=ZERO; digit3<=NINE; end
      16'd9020: begin digit0<=ZERO; digit1<=TWO; digit2<=ZERO; digit3<=NINE; end
      16'd9021: begin digit0<=ONE; digit1<=TWO; digit2<=ZERO; digit3<=NINE; end
      16'd9022: begin digit0<=TWO; digit1<=TWO; digit2<=ZERO; digit3<=NINE; end
      16'd9023: begin digit0<=THREE; digit1<=TWO; digit2<=ZERO; digit3<=NINE; end
      16'd9024: begin digit0<=FOUR; digit1<=TWO; digit2<=ZERO; digit3<=NINE; end
      16'd9025: begin digit0<=FIVE; digit1<=TWO; digit2<=ZERO; digit3<=NINE; end
      16'd9026: begin digit0<=SIX; digit1<=TWO; digit2<=ZERO; digit3<=NINE; end
      16'd9027: begin digit0<=SEVEN; digit1<=TWO; digit2<=ZERO; digit3<=NINE; end
      16'd9028: begin digit0<=EIGHT; digit1<=TWO; digit2<=ZERO; digit3<=NINE; end
      16'd9029: begin digit0<=NINE; digit1<=TWO; digit2<=ZERO; digit3<=NINE; end
      16'd9030: begin digit0<=ZERO; digit1<=THREE; digit2<=ZERO; digit3<=NINE; end
      16'd9031: begin digit0<=ONE; digit1<=THREE; digit2<=ZERO; digit3<=NINE; end
      16'd9032: begin digit0<=TWO; digit1<=THREE; digit2<=ZERO; digit3<=NINE; end
      16'd9033: begin digit0<=THREE; digit1<=THREE; digit2<=ZERO; digit3<=NINE; end
      16'd9034: begin digit0<=FOUR; digit1<=THREE; digit2<=ZERO; digit3<=NINE; end
      16'd9035: begin digit0<=FIVE; digit1<=THREE; digit2<=ZERO; digit3<=NINE; end
      16'd9036: begin digit0<=SIX; digit1<=THREE; digit2<=ZERO; digit3<=NINE; end
      16'd9037: begin digit0<=SEVEN; digit1<=THREE; digit2<=ZERO; digit3<=NINE; end
      16'd9038: begin digit0<=EIGHT; digit1<=THREE; digit2<=ZERO; digit3<=NINE; end
      16'd9039: begin digit0<=NINE; digit1<=THREE; digit2<=ZERO; digit3<=NINE; end
      16'd9040: begin digit0<=ZERO; digit1<=FOUR; digit2<=ZERO; digit3<=NINE; end
      16'd9041: begin digit0<=ONE; digit1<=FOUR; digit2<=ZERO; digit3<=NINE; end
      16'd9042: begin digit0<=TWO; digit1<=FOUR; digit2<=ZERO; digit3<=NINE; end
      16'd9043: begin digit0<=THREE; digit1<=FOUR; digit2<=ZERO; digit3<=NINE; end
      16'd9044: begin digit0<=FOUR; digit1<=FOUR; digit2<=ZERO; digit3<=NINE; end
      16'd9045: begin digit0<=FIVE; digit1<=FOUR; digit2<=ZERO; digit3<=NINE; end
      16'd9046: begin digit0<=SIX; digit1<=FOUR; digit2<=ZERO; digit3<=NINE; end
      16'd9047: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ZERO; digit3<=NINE; end
      16'd9048: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ZERO; digit3<=NINE; end
      16'd9049: begin digit0<=NINE; digit1<=FOUR; digit2<=ZERO; digit3<=NINE; end
      16'd9050: begin digit0<=ZERO; digit1<=FIVE; digit2<=ZERO; digit3<=NINE; end
      16'd9051: begin digit0<=ONE; digit1<=FIVE; digit2<=ZERO; digit3<=NINE; end
      16'd9052: begin digit0<=TWO; digit1<=FIVE; digit2<=ZERO; digit3<=NINE; end
      16'd9053: begin digit0<=THREE; digit1<=FIVE; digit2<=ZERO; digit3<=NINE; end
      16'd9054: begin digit0<=FOUR; digit1<=FIVE; digit2<=ZERO; digit3<=NINE; end
      16'd9055: begin digit0<=FIVE; digit1<=FIVE; digit2<=ZERO; digit3<=NINE; end
      16'd9056: begin digit0<=SIX; digit1<=FIVE; digit2<=ZERO; digit3<=NINE; end
      16'd9057: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ZERO; digit3<=NINE; end
      16'd9058: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ZERO; digit3<=NINE; end
      16'd9059: begin digit0<=NINE; digit1<=FIVE; digit2<=ZERO; digit3<=NINE; end
      16'd9060: begin digit0<=ZERO; digit1<=SIX; digit2<=ZERO; digit3<=NINE; end
      16'd9061: begin digit0<=ONE; digit1<=SIX; digit2<=ZERO; digit3<=NINE; end
      16'd9062: begin digit0<=TWO; digit1<=SIX; digit2<=ZERO; digit3<=NINE; end
      16'd9063: begin digit0<=THREE; digit1<=SIX; digit2<=ZERO; digit3<=NINE; end
      16'd9064: begin digit0<=FOUR; digit1<=SIX; digit2<=ZERO; digit3<=NINE; end
      16'd9065: begin digit0<=FIVE; digit1<=SIX; digit2<=ZERO; digit3<=NINE; end
      16'd9066: begin digit0<=SIX; digit1<=SIX; digit2<=ZERO; digit3<=NINE; end
      16'd9067: begin digit0<=SEVEN; digit1<=SIX; digit2<=ZERO; digit3<=NINE; end
      16'd9068: begin digit0<=EIGHT; digit1<=SIX; digit2<=ZERO; digit3<=NINE; end
      16'd9069: begin digit0<=NINE; digit1<=SIX; digit2<=ZERO; digit3<=NINE; end
      16'd9070: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ZERO; digit3<=NINE; end
      16'd9071: begin digit0<=ONE; digit1<=SEVEN; digit2<=ZERO; digit3<=NINE; end
      16'd9072: begin digit0<=TWO; digit1<=SEVEN; digit2<=ZERO; digit3<=NINE; end
      16'd9073: begin digit0<=THREE; digit1<=SEVEN; digit2<=ZERO; digit3<=NINE; end
      16'd9074: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ZERO; digit3<=NINE; end
      16'd9075: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ZERO; digit3<=NINE; end
      16'd9076: begin digit0<=SIX; digit1<=SEVEN; digit2<=ZERO; digit3<=NINE; end
      16'd9077: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ZERO; digit3<=NINE; end
      16'd9078: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ZERO; digit3<=NINE; end
      16'd9079: begin digit0<=NINE; digit1<=SEVEN; digit2<=ZERO; digit3<=NINE; end
      16'd9080: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ZERO; digit3<=NINE; end
      16'd9081: begin digit0<=ONE; digit1<=EIGHT; digit2<=ZERO; digit3<=NINE; end
      16'd9082: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ZERO; digit3<=NINE; end
      16'd9083: begin digit0<=THREE; digit1<=EIGHT; digit2<=ZERO; digit3<=NINE; end
      16'd9084: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ZERO; digit3<=NINE; end
      16'd9085: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ZERO; digit3<=NINE; end
      16'd9086: begin digit0<=SIX; digit1<=EIGHT; digit2<=ZERO; digit3<=NINE; end
      16'd9087: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ZERO; digit3<=NINE; end
      16'd9088: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ZERO; digit3<=NINE; end
      16'd9089: begin digit0<=NINE; digit1<=EIGHT; digit2<=ZERO; digit3<=NINE; end
      16'd9090: begin digit0<=ZERO; digit1<=NINE; digit2<=ZERO; digit3<=NINE; end
      16'd9091: begin digit0<=ONE; digit1<=NINE; digit2<=ZERO; digit3<=NINE; end
      16'd9092: begin digit0<=ZERO; digit1<=NINE; digit2<=ZERO; digit3<=NINE; end
      16'd9093: begin digit0<=THREE; digit1<=NINE; digit2<=ZERO; digit3<=NINE; end
      16'd9094: begin digit0<=FOUR; digit1<=NINE; digit2<=ZERO; digit3<=NINE; end
      16'd9095: begin digit0<=FIVE; digit1<=NINE; digit2<=ZERO; digit3<=NINE; end
      16'd9096: begin digit0<=SIX; digit1<=NINE; digit2<=ZERO; digit3<=NINE; end
      16'd9097: begin digit0<=SEVEN; digit1<=NINE; digit2<=ZERO; digit3<=NINE; end
      16'd9098: begin digit0<=EIGHT; digit1<=NINE; digit2<=ZERO; digit3<=NINE; end
      16'd9099: begin digit0<=NINE; digit1<=NINE; digit2<=ZERO; digit3<=NINE; end
	  16'd9100: begin digit0<=ZERO; digit1<=ZERO; digit2<=ONE; digit3<=NINE; end
      16'd9101: begin digit0<=ONE; digit1<=ZERO; digit2<=ONE; digit3<=NINE; end
      16'd9102: begin digit0<=TWO; digit1<=ZERO; digit2<=ONE; digit3<=NINE; end
      16'd9103: begin digit0<=THREE; digit1<=ZERO; digit2<=ONE; digit3<=NINE; end
      16'd9104: begin digit0<=FOUR; digit1<=ZERO; digit2<=ONE; digit3<=NINE; end
      16'd9105: begin digit0<=FIVE; digit1<=ZERO; digit2<=ONE; digit3<=NINE; end
      16'd9106: begin digit0<=SIX; digit1<=ZERO; digit2<=ONE; digit3<=NINE; end
      16'd9107: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ONE; digit3<=NINE; end
      16'd9108: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ONE; digit3<=NINE; end
      16'd9109: begin digit0<=NINE; digit1<=ZERO; digit2<=ONE; digit3<=NINE; end
      16'd9110: begin digit0<=ZERO; digit1<=ONE; digit2<=ONE; digit3<=NINE; end
      16'd9111: begin digit0<=ONE; digit1<=ONE; digit2<=ONE; digit3<=NINE; end
      16'd9112: begin digit0<=TWO; digit1<=ONE; digit2<=ONE; digit3<=NINE; end
      16'd9113: begin digit0<=THREE; digit1<=ONE; digit2<=ONE; digit3<=NINE; end
      16'd9114: begin digit0<=FOUR; digit1<=ONE; digit2<=ONE; digit3<=NINE; end
      16'd9115: begin digit0<=FIVE; digit1<=ONE; digit2<=ONE; digit3<=NINE; end
      16'd9116: begin digit0<=SIX; digit1<=ONE; digit2<=ONE; digit3<=NINE; end
      16'd9117: begin digit0<=SEVEN; digit1<=ONE; digit2<=ONE; digit3<=NINE; end
      16'd9118: begin digit0<=EIGHT; digit1<=ONE; digit2<=ONE; digit3<=NINE; end
      16'd9119: begin digit0<=NINE; digit1<=ONE; digit2<=ONE; digit3<=NINE; end
      16'd9120: begin digit0<=ZERO; digit1<=TWO; digit2<=ONE; digit3<=NINE; end
      16'd9121: begin digit0<=ONE; digit1<=TWO; digit2<=ONE; digit3<=NINE; end
      16'd9122: begin digit0<=TWO; digit1<=TWO; digit2<=ONE; digit3<=NINE; end
      16'd9123: begin digit0<=THREE; digit1<=TWO; digit2<=ONE; digit3<=NINE; end
      16'd9124: begin digit0<=FOUR; digit1<=TWO; digit2<=ONE; digit3<=NINE; end
      16'd9125: begin digit0<=FIVE; digit1<=TWO; digit2<=ONE; digit3<=NINE; end
      16'd9126: begin digit0<=SIX; digit1<=TWO; digit2<=ONE; digit3<=NINE; end
      16'd9127: begin digit0<=SEVEN; digit1<=TWO; digit2<=ONE; digit3<=NINE; end
      16'd9128: begin digit0<=EIGHT; digit1<=TWO; digit2<=ONE; digit3<=NINE; end
      16'd9129: begin digit0<=NINE; digit1<=TWO; digit2<=ONE; digit3<=NINE; end
      16'd9130: begin digit0<=ZERO; digit1<=THREE; digit2<=ONE; digit3<=NINE; end
      16'd9131: begin digit0<=ONE; digit1<=THREE; digit2<=ONE; digit3<=NINE; end
      16'd9132: begin digit0<=TWO; digit1<=THREE; digit2<=ONE; digit3<=NINE; end
      16'd9133: begin digit0<=THREE; digit1<=THREE; digit2<=ONE; digit3<=NINE; end
      16'd9134: begin digit0<=FOUR; digit1<=THREE; digit2<=ONE; digit3<=NINE; end
      16'd9135: begin digit0<=FIVE; digit1<=THREE; digit2<=ONE; digit3<=NINE; end
      16'd9136: begin digit0<=SIX; digit1<=THREE; digit2<=ONE; digit3<=NINE; end
      16'd9137: begin digit0<=SEVEN; digit1<=THREE; digit2<=ONE; digit3<=NINE; end
      16'd9138: begin digit0<=EIGHT; digit1<=THREE; digit2<=ONE; digit3<=NINE; end
      16'd9139: begin digit0<=NINE; digit1<=THREE; digit2<=ONE; digit3<=NINE; end
      16'd9140: begin digit0<=ZERO; digit1<=FOUR; digit2<=ONE; digit3<=NINE; end
      16'd9141: begin digit0<=ONE; digit1<=FOUR; digit2<=ONE; digit3<=NINE; end
      16'd9142: begin digit0<=TWO; digit1<=FOUR; digit2<=ONE; digit3<=NINE; end
      16'd9143: begin digit0<=THREE; digit1<=FOUR; digit2<=ONE; digit3<=NINE; end
      16'd9144: begin digit0<=FOUR; digit1<=FOUR; digit2<=ONE; digit3<=NINE; end
      16'd9145: begin digit0<=FIVE; digit1<=FOUR; digit2<=ONE; digit3<=NINE; end
      16'd9146: begin digit0<=SIX; digit1<=FOUR; digit2<=ONE; digit3<=NINE; end
      16'd9147: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ONE; digit3<=NINE; end
      16'd9148: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ONE; digit3<=NINE; end
      16'd9149: begin digit0<=NINE; digit1<=FOUR; digit2<=ONE; digit3<=NINE; end
      16'd9150: begin digit0<=ZERO; digit1<=FIVE; digit2<=ONE; digit3<=NINE; end
      16'd9151: begin digit0<=ONE; digit1<=FIVE; digit2<=ONE; digit3<=NINE; end
      16'd9152: begin digit0<=TWO; digit1<=FIVE; digit2<=ONE; digit3<=NINE; end
      16'd9153: begin digit0<=THREE; digit1<=FIVE; digit2<=ONE; digit3<=NINE; end
      16'd9154: begin digit0<=FOUR; digit1<=FIVE; digit2<=ONE; digit3<=NINE; end
      16'd9155: begin digit0<=FIVE; digit1<=FIVE; digit2<=ONE; digit3<=NINE; end
      16'd9156: begin digit0<=SIX; digit1<=FIVE; digit2<=ONE; digit3<=NINE; end
      16'd9157: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ONE; digit3<=NINE; end
      16'd9158: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ONE; digit3<=NINE; end
      16'd9159: begin digit0<=NINE; digit1<=FIVE; digit2<=ONE; digit3<=NINE; end
      16'd9160: begin digit0<=ZERO; digit1<=SIX; digit2<=ONE; digit3<=NINE; end
      16'd9161: begin digit0<=ONE; digit1<=SIX; digit2<=ONE; digit3<=NINE; end
      16'd9162: begin digit0<=TWO; digit1<=SIX; digit2<=ONE; digit3<=NINE; end
      16'd9163: begin digit0<=THREE; digit1<=SIX; digit2<=ONE; digit3<=NINE; end
      16'd9164: begin digit0<=FOUR; digit1<=SIX; digit2<=ONE; digit3<=NINE; end
      16'd9165: begin digit0<=FIVE; digit1<=SIX; digit2<=ONE; digit3<=NINE; end
      16'd9166: begin digit0<=SIX; digit1<=SIX; digit2<=ONE; digit3<=NINE; end
      16'd9167: begin digit0<=SEVEN; digit1<=SIX; digit2<=ONE; digit3<=NINE; end
      16'd9168: begin digit0<=EIGHT; digit1<=SIX; digit2<=ONE; digit3<=NINE; end
      16'd9169: begin digit0<=NINE; digit1<=SIX; digit2<=ONE; digit3<=NINE; end
      16'd9170: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ONE; digit3<=NINE; end
      16'd9171: begin digit0<=ONE; digit1<=SEVEN; digit2<=ONE; digit3<=NINE; end
      16'd9172: begin digit0<=TWO; digit1<=SEVEN; digit2<=ONE; digit3<=NINE; end
      16'd9173: begin digit0<=THREE; digit1<=SEVEN; digit2<=ONE; digit3<=NINE; end
      16'd9174: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ONE; digit3<=NINE; end
      16'd9175: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ONE; digit3<=NINE; end
      16'd9176: begin digit0<=SIX; digit1<=SEVEN; digit2<=ONE; digit3<=NINE; end
      16'd9177: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ONE; digit3<=NINE; end
      16'd9178: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ONE; digit3<=NINE; end
      16'd9179: begin digit0<=NINE; digit1<=SEVEN; digit2<=ONE; digit3<=NINE; end
      16'd9180: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=NINE; end
      16'd9181: begin digit0<=ONE; digit1<=EIGHT; digit2<=ONE; digit3<=NINE; end
      16'd9182: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=NINE; end
      16'd9183: begin digit0<=THREE; digit1<=EIGHT; digit2<=ONE; digit3<=NINE; end
      16'd9184: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ONE; digit3<=NINE; end
      16'd9185: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ONE; digit3<=NINE; end
      16'd9186: begin digit0<=SIX; digit1<=EIGHT; digit2<=ONE; digit3<=NINE; end
      16'd9187: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ONE; digit3<=NINE; end
      16'd9188: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ONE; digit3<=NINE; end
      16'd9189: begin digit0<=NINE; digit1<=EIGHT; digit2<=ONE; digit3<=NINE; end
      16'd9190: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=NINE; end
      16'd9191: begin digit0<=ONE; digit1<=NINE; digit2<=ONE; digit3<=NINE; end
      16'd9192: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=NINE; end
      16'd9193: begin digit0<=THREE; digit1<=NINE; digit2<=ONE; digit3<=NINE; end
      16'd9194: begin digit0<=FOUR; digit1<=NINE; digit2<=ONE; digit3<=NINE; end
      16'd9195: begin digit0<=FIVE; digit1<=NINE; digit2<=ONE; digit3<=NINE; end
      16'd9196: begin digit0<=SIX; digit1<=NINE; digit2<=ONE; digit3<=NINE; end
      16'd9197: begin digit0<=SEVEN; digit1<=NINE; digit2<=ONE; digit3<=NINE; end
      16'd9198: begin digit0<=EIGHT; digit1<=NINE; digit2<=ONE; digit3<=NINE; end
      16'd9199: begin digit0<=NINE; digit1<=NINE; digit2<=ONE; digit3<=NINE; end
	  16'd9200: begin digit0<=ZERO; digit1<=ZERO; digit2<=TWO; digit3<=NINE; end
      16'd9201: begin digit0<=ONE; digit1<=ZERO; digit2<=TWO; digit3<=NINE; end
      16'd9202: begin digit0<=TWO; digit1<=ZERO; digit2<=TWO; digit3<=NINE; end
      16'd9203: begin digit0<=THREE; digit1<=ZERO; digit2<=TWO; digit3<=NINE; end
      16'd9204: begin digit0<=FOUR; digit1<=ZERO; digit2<=TWO; digit3<=NINE; end
      16'd9205: begin digit0<=FIVE; digit1<=ZERO; digit2<=TWO; digit3<=NINE; end
      16'd9206: begin digit0<=SIX; digit1<=ZERO; digit2<=TWO; digit3<=NINE; end
      16'd9207: begin digit0<=SEVEN; digit1<=ZERO; digit2<=TWO; digit3<=NINE; end
      16'd9208: begin digit0<=EIGHT; digit1<=ZERO; digit2<=TWO; digit3<=NINE; end
      16'd9209: begin digit0<=NINE; digit1<=ZERO; digit2<=TWO; digit3<=NINE; end
      16'd9210: begin digit0<=ZERO; digit1<=ONE; digit2<=TWO; digit3<=NINE; end
      16'd9211: begin digit0<=ONE; digit1<=ONE; digit2<=TWO; digit3<=NINE; end
      16'd9212: begin digit0<=TWO; digit1<=ONE; digit2<=TWO; digit3<=NINE; end
      16'd9213: begin digit0<=THREE; digit1<=ONE; digit2<=TWO; digit3<=NINE; end
      16'd9214: begin digit0<=FOUR; digit1<=ONE; digit2<=TWO; digit3<=NINE; end
      16'd9215: begin digit0<=FIVE; digit1<=ONE; digit2<=TWO; digit3<=NINE; end
      16'd9216: begin digit0<=SIX; digit1<=ONE; digit2<=TWO; digit3<=NINE; end
      16'd9217: begin digit0<=SEVEN; digit1<=ONE; digit2<=TWO; digit3<=NINE; end
      16'd9218: begin digit0<=EIGHT; digit1<=ONE; digit2<=TWO; digit3<=NINE; end
      16'd9219: begin digit0<=NINE; digit1<=ONE; digit2<=TWO; digit3<=NINE; end
      16'd9220: begin digit0<=ZERO; digit1<=TWO; digit2<=TWO; digit3<=NINE; end
      16'd9221: begin digit0<=ONE; digit1<=TWO; digit2<=TWO; digit3<=NINE; end
      16'd9222: begin digit0<=TWO; digit1<=TWO; digit2<=TWO; digit3<=NINE; end
      16'd9223: begin digit0<=THREE; digit1<=TWO; digit2<=TWO; digit3<=NINE; end
      16'd9224: begin digit0<=FOUR; digit1<=TWO; digit2<=TWO; digit3<=NINE; end
      16'd9225: begin digit0<=FIVE; digit1<=TWO; digit2<=TWO; digit3<=NINE; end
      16'd9226: begin digit0<=SIX; digit1<=TWO; digit2<=TWO; digit3<=NINE; end
      16'd9227: begin digit0<=SEVEN; digit1<=TWO; digit2<=TWO; digit3<=NINE; end
      16'd9228: begin digit0<=EIGHT; digit1<=TWO; digit2<=TWO; digit3<=NINE; end
      16'd9229: begin digit0<=NINE; digit1<=TWO; digit2<=TWO; digit3<=NINE; end
      16'd9230: begin digit0<=ZERO; digit1<=THREE; digit2<=TWO; digit3<=NINE; end
      16'd9231: begin digit0<=ONE; digit1<=THREE; digit2<=TWO; digit3<=NINE; end
      16'd9232: begin digit0<=TWO; digit1<=THREE; digit2<=TWO; digit3<=NINE; end
      16'd9233: begin digit0<=THREE; digit1<=THREE; digit2<=TWO; digit3<=NINE; end
      16'd9234: begin digit0<=FOUR; digit1<=THREE; digit2<=TWO; digit3<=NINE; end
      16'd9235: begin digit0<=FIVE; digit1<=THREE; digit2<=TWO; digit3<=NINE; end
      16'd9236: begin digit0<=SIX; digit1<=THREE; digit2<=TWO; digit3<=NINE; end
      16'd9237: begin digit0<=SEVEN; digit1<=THREE; digit2<=TWO; digit3<=NINE; end
      16'd9238: begin digit0<=EIGHT; digit1<=THREE; digit2<=TWO; digit3<=NINE; end
      16'd9239: begin digit0<=NINE; digit1<=THREE; digit2<=TWO; digit3<=NINE; end
      16'd9240: begin digit0<=ZERO; digit1<=FOUR; digit2<=TWO; digit3<=NINE; end
      16'd9241: begin digit0<=ONE; digit1<=FOUR; digit2<=TWO; digit3<=NINE; end
      16'd9242: begin digit0<=TWO; digit1<=FOUR; digit2<=TWO; digit3<=NINE; end
      16'd9243: begin digit0<=THREE; digit1<=FOUR; digit2<=TWO; digit3<=NINE; end
      16'd9244: begin digit0<=FOUR; digit1<=FOUR; digit2<=TWO; digit3<=NINE; end
      16'd9245: begin digit0<=FIVE; digit1<=FOUR; digit2<=TWO; digit3<=NINE; end
      16'd9246: begin digit0<=SIX; digit1<=FOUR; digit2<=TWO; digit3<=NINE; end
      16'd9247: begin digit0<=SEVEN; digit1<=FOUR; digit2<=TWO; digit3<=NINE; end
      16'd9248: begin digit0<=EIGHT; digit1<=FOUR; digit2<=TWO; digit3<=NINE; end
      16'd9249: begin digit0<=NINE; digit1<=FOUR; digit2<=TWO; digit3<=NINE; end
      16'd9250: begin digit0<=ZERO; digit1<=FIVE; digit2<=TWO; digit3<=NINE; end
      16'd9251: begin digit0<=ONE; digit1<=FIVE; digit2<=TWO; digit3<=NINE; end
      16'd9252: begin digit0<=TWO; digit1<=FIVE; digit2<=TWO; digit3<=NINE; end
      16'd9253: begin digit0<=THREE; digit1<=FIVE; digit2<=TWO; digit3<=NINE; end
      16'd9254: begin digit0<=FOUR; digit1<=FIVE; digit2<=TWO; digit3<=NINE; end
      16'd9255: begin digit0<=FIVE; digit1<=FIVE; digit2<=TWO; digit3<=NINE; end
      16'd9256: begin digit0<=SIX; digit1<=FIVE; digit2<=TWO; digit3<=NINE; end
      16'd9257: begin digit0<=SEVEN; digit1<=FIVE; digit2<=TWO; digit3<=NINE; end
      16'd9258: begin digit0<=EIGHT; digit1<=FIVE; digit2<=TWO; digit3<=NINE; end
      16'd9259: begin digit0<=NINE; digit1<=FIVE; digit2<=TWO; digit3<=NINE; end
      16'd9260: begin digit0<=ZERO; digit1<=SIX; digit2<=TWO; digit3<=NINE; end
      16'd9261: begin digit0<=ONE; digit1<=SIX; digit2<=TWO; digit3<=NINE; end
      16'd9262: begin digit0<=TWO; digit1<=SIX; digit2<=TWO; digit3<=NINE; end
      16'd9263: begin digit0<=THREE; digit1<=SIX; digit2<=TWO; digit3<=NINE; end
      16'd9264: begin digit0<=FOUR; digit1<=SIX; digit2<=TWO; digit3<=NINE; end
      16'd9265: begin digit0<=FIVE; digit1<=SIX; digit2<=TWO; digit3<=NINE; end
      16'd9266: begin digit0<=SIX; digit1<=SIX; digit2<=TWO; digit3<=NINE; end
      16'd9267: begin digit0<=SEVEN; digit1<=SIX; digit2<=TWO; digit3<=NINE; end
      16'd9268: begin digit0<=EIGHT; digit1<=SIX; digit2<=TWO; digit3<=NINE; end
      16'd9269: begin digit0<=NINE; digit1<=SIX; digit2<=TWO; digit3<=NINE; end
      16'd9270: begin digit0<=ZERO; digit1<=SEVEN; digit2<=TWO; digit3<=NINE; end
      16'd9271: begin digit0<=ONE; digit1<=SEVEN; digit2<=TWO; digit3<=NINE; end
      16'd9272: begin digit0<=TWO; digit1<=SEVEN; digit2<=TWO; digit3<=NINE; end
      16'd9273: begin digit0<=THREE; digit1<=SEVEN; digit2<=TWO; digit3<=NINE; end
      16'd9274: begin digit0<=FOUR; digit1<=SEVEN; digit2<=TWO; digit3<=NINE; end
      16'd9275: begin digit0<=FIVE; digit1<=SEVEN; digit2<=TWO; digit3<=NINE; end
      16'd9276: begin digit0<=SIX; digit1<=SEVEN; digit2<=TWO; digit3<=NINE; end
      16'd9277: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=TWO; digit3<=NINE; end
      16'd9278: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=TWO; digit3<=NINE; end
      16'd9279: begin digit0<=NINE; digit1<=SEVEN; digit2<=TWO; digit3<=NINE; end
      16'd9280: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=NINE; end
      16'd9281: begin digit0<=ONE; digit1<=EIGHT; digit2<=TWO; digit3<=NINE; end
      16'd9282: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=NINE; end
      16'd9283: begin digit0<=THREE; digit1<=EIGHT; digit2<=TWO; digit3<=NINE; end
      16'd9284: begin digit0<=FOUR; digit1<=EIGHT; digit2<=TWO; digit3<=NINE; end
      16'd9285: begin digit0<=FIVE; digit1<=EIGHT; digit2<=TWO; digit3<=NINE; end
      16'd9286: begin digit0<=SIX; digit1<=EIGHT; digit2<=TWO; digit3<=NINE; end
      16'd9287: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=TWO; digit3<=NINE; end
      16'd9288: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=TWO; digit3<=NINE; end
      16'd9289: begin digit0<=NINE; digit1<=EIGHT; digit2<=TWO; digit3<=NINE; end
      16'd9290: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=NINE; end
      16'd9291: begin digit0<=ONE; digit1<=NINE; digit2<=TWO; digit3<=NINE; end
      16'd9292: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=NINE; end
      16'd9293: begin digit0<=THREE; digit1<=NINE; digit2<=TWO; digit3<=NINE; end
      16'd9294: begin digit0<=FOUR; digit1<=NINE; digit2<=TWO; digit3<=NINE; end
      16'd9295: begin digit0<=FIVE; digit1<=NINE; digit2<=TWO; digit3<=NINE; end
      16'd9296: begin digit0<=SIX; digit1<=NINE; digit2<=TWO; digit3<=NINE; end
      16'd9297: begin digit0<=SEVEN; digit1<=NINE; digit2<=TWO; digit3<=NINE; end
      16'd9298: begin digit0<=EIGHT; digit1<=NINE; digit2<=TWO; digit3<=NINE; end
      16'd9299: begin digit0<=NINE; digit1<=NINE; digit2<=TWO; digit3<=NINE; end
	  16'd9300: begin digit0<=ZERO; digit1<=ZERO; digit2<=THREE; digit3<=NINE; end
      16'd9301: begin digit0<=ONE; digit1<=ZERO; digit2<=THREE; digit3<=NINE; end
      16'd9302: begin digit0<=TWO; digit1<=ZERO; digit2<=THREE; digit3<=NINE; end
      16'd9303: begin digit0<=THREE; digit1<=ZERO; digit2<=THREE; digit3<=NINE; end
      16'd9304: begin digit0<=FOUR; digit1<=ZERO; digit2<=THREE; digit3<=NINE; end
      16'd9305: begin digit0<=FIVE; digit1<=ZERO; digit2<=THREE; digit3<=NINE; end
      16'd9306: begin digit0<=SIX; digit1<=ZERO; digit2<=THREE; digit3<=NINE; end
      16'd9307: begin digit0<=SEVEN; digit1<=ZERO; digit2<=THREE; digit3<=NINE; end
      16'd9308: begin digit0<=EIGHT; digit1<=ZERO; digit2<=THREE; digit3<=NINE; end
      16'd9309: begin digit0<=NINE; digit1<=ZERO; digit2<=THREE; digit3<=NINE; end
      16'd9310: begin digit0<=ZERO; digit1<=ONE; digit2<=THREE; digit3<=NINE; end
      16'd9311: begin digit0<=ONE; digit1<=ONE; digit2<=THREE; digit3<=NINE; end
      16'd9312: begin digit0<=TWO; digit1<=ONE; digit2<=THREE; digit3<=NINE; end
      16'd9313: begin digit0<=THREE; digit1<=ONE; digit2<=THREE; digit3<=NINE; end
      16'd9314: begin digit0<=FOUR; digit1<=ONE; digit2<=THREE; digit3<=NINE; end
      16'd9315: begin digit0<=FIVE; digit1<=ONE; digit2<=THREE; digit3<=NINE; end
      16'd9316: begin digit0<=SIX; digit1<=ONE; digit2<=THREE; digit3<=NINE; end
      16'd9317: begin digit0<=SEVEN; digit1<=ONE; digit2<=THREE; digit3<=NINE; end
      16'd9318: begin digit0<=EIGHT; digit1<=ONE; digit2<=THREE; digit3<=NINE; end
      16'd9319: begin digit0<=NINE; digit1<=ONE; digit2<=THREE; digit3<=NINE; end
      16'd9320: begin digit0<=ZERO; digit1<=TWO; digit2<=THREE; digit3<=NINE; end
      16'd9321: begin digit0<=ONE; digit1<=TWO; digit2<=THREE; digit3<=NINE; end
      16'd9322: begin digit0<=TWO; digit1<=TWO; digit2<=THREE; digit3<=NINE; end
      16'd9323: begin digit0<=THREE; digit1<=TWO; digit2<=THREE; digit3<=NINE; end
      16'd9324: begin digit0<=FOUR; digit1<=TWO; digit2<=THREE; digit3<=NINE; end
      16'd9325: begin digit0<=FIVE; digit1<=TWO; digit2<=THREE; digit3<=NINE; end
      16'd9326: begin digit0<=SIX; digit1<=TWO; digit2<=THREE; digit3<=NINE; end
      16'd9327: begin digit0<=SEVEN; digit1<=TWO; digit2<=THREE; digit3<=NINE; end
      16'd9328: begin digit0<=EIGHT; digit1<=TWO; digit2<=THREE; digit3<=NINE; end
      16'd9329: begin digit0<=NINE; digit1<=TWO; digit2<=THREE; digit3<=NINE; end
      16'd9330: begin digit0<=ZERO; digit1<=THREE; digit2<=THREE; digit3<=NINE; end
      16'd9331: begin digit0<=ONE; digit1<=THREE; digit2<=THREE; digit3<=NINE; end
      16'd9332: begin digit0<=TWO; digit1<=THREE; digit2<=THREE; digit3<=NINE; end
      16'd9333: begin digit0<=THREE; digit1<=THREE; digit2<=THREE; digit3<=NINE; end
      16'd9334: begin digit0<=FOUR; digit1<=THREE; digit2<=THREE; digit3<=NINE; end
      16'd9335: begin digit0<=FIVE; digit1<=THREE; digit2<=THREE; digit3<=NINE; end
      16'd9336: begin digit0<=SIX; digit1<=THREE; digit2<=THREE; digit3<=NINE; end
      16'd9337: begin digit0<=SEVEN; digit1<=THREE; digit2<=THREE; digit3<=NINE; end
      16'd9338: begin digit0<=EIGHT; digit1<=THREE; digit2<=THREE; digit3<=NINE; end
      16'd9339: begin digit0<=NINE; digit1<=THREE; digit2<=THREE; digit3<=NINE; end
      16'd9340: begin digit0<=ZERO; digit1<=FOUR; digit2<=THREE; digit3<=NINE; end
      16'd9341: begin digit0<=ONE; digit1<=FOUR; digit2<=THREE; digit3<=NINE; end
      16'd9342: begin digit0<=TWO; digit1<=FOUR; digit2<=THREE; digit3<=NINE; end
      16'd9343: begin digit0<=THREE; digit1<=FOUR; digit2<=THREE; digit3<=NINE; end
      16'd9344: begin digit0<=FOUR; digit1<=FOUR; digit2<=THREE; digit3<=NINE; end
      16'd9345: begin digit0<=FIVE; digit1<=FOUR; digit2<=THREE; digit3<=NINE; end
      16'd9346: begin digit0<=SIX; digit1<=FOUR; digit2<=THREE; digit3<=NINE; end
      16'd9347: begin digit0<=SEVEN; digit1<=FOUR; digit2<=THREE; digit3<=NINE; end
      16'd9348: begin digit0<=EIGHT; digit1<=FOUR; digit2<=THREE; digit3<=NINE; end
      16'd9349: begin digit0<=NINE; digit1<=FOUR; digit2<=THREE; digit3<=NINE; end
      16'd9350: begin digit0<=ZERO; digit1<=FIVE; digit2<=THREE; digit3<=NINE; end
      16'd9351: begin digit0<=ONE; digit1<=FIVE; digit2<=THREE; digit3<=NINE; end
      16'd9352: begin digit0<=TWO; digit1<=FIVE; digit2<=THREE; digit3<=NINE; end
      16'd9353: begin digit0<=THREE; digit1<=FIVE; digit2<=THREE; digit3<=NINE; end
      16'd9354: begin digit0<=FOUR; digit1<=FIVE; digit2<=THREE; digit3<=NINE; end
      16'd9355: begin digit0<=FIVE; digit1<=FIVE; digit2<=THREE; digit3<=NINE; end
      16'd9356: begin digit0<=SIX; digit1<=FIVE; digit2<=THREE; digit3<=NINE; end
      16'd9357: begin digit0<=SEVEN; digit1<=FIVE; digit2<=THREE; digit3<=NINE; end
      16'd9358: begin digit0<=EIGHT; digit1<=FIVE; digit2<=THREE; digit3<=NINE; end
      16'd9359: begin digit0<=NINE; digit1<=FIVE; digit2<=THREE; digit3<=NINE; end
      16'd9360: begin digit0<=ZERO; digit1<=SIX; digit2<=THREE; digit3<=NINE; end
      16'd9361: begin digit0<=ONE; digit1<=SIX; digit2<=THREE; digit3<=NINE; end
      16'd9362: begin digit0<=TWO; digit1<=SIX; digit2<=THREE; digit3<=NINE; end
      16'd9363: begin digit0<=THREE; digit1<=SIX; digit2<=THREE; digit3<=NINE; end
      16'd9364: begin digit0<=FOUR; digit1<=SIX; digit2<=THREE; digit3<=NINE; end
      16'd9365: begin digit0<=FIVE; digit1<=SIX; digit2<=THREE; digit3<=NINE; end
      16'd9366: begin digit0<=SIX; digit1<=SIX; digit2<=THREE; digit3<=NINE; end
      16'd9367: begin digit0<=SEVEN; digit1<=SIX; digit2<=THREE; digit3<=NINE; end
      16'd9368: begin digit0<=EIGHT; digit1<=SIX; digit2<=THREE; digit3<=NINE; end
      16'd9369: begin digit0<=NINE; digit1<=SIX; digit2<=THREE; digit3<=NINE; end
      16'd9370: begin digit0<=ZERO; digit1<=SEVEN; digit2<=THREE; digit3<=NINE; end
      16'd9371: begin digit0<=ONE; digit1<=SEVEN; digit2<=THREE; digit3<=NINE; end
      16'd9372: begin digit0<=TWO; digit1<=SEVEN; digit2<=THREE; digit3<=NINE; end
      16'd9373: begin digit0<=THREE; digit1<=SEVEN; digit2<=THREE; digit3<=NINE; end
      16'd9374: begin digit0<=FOUR; digit1<=SEVEN; digit2<=THREE; digit3<=NINE; end
      16'd9375: begin digit0<=FIVE; digit1<=SEVEN; digit2<=THREE; digit3<=NINE; end
      16'd9376: begin digit0<=SIX; digit1<=SEVEN; digit2<=THREE; digit3<=NINE; end
      16'd9377: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=THREE; digit3<=NINE; end
      16'd9378: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=THREE; digit3<=NINE; end
      16'd9379: begin digit0<=NINE; digit1<=SEVEN; digit2<=THREE; digit3<=NINE; end
      16'd9380: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=NINE; end
      16'd9381: begin digit0<=ONE; digit1<=EIGHT; digit2<=THREE; digit3<=NINE; end
      16'd9382: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=NINE; end
      16'd9383: begin digit0<=THREE; digit1<=EIGHT; digit2<=THREE; digit3<=NINE; end
      16'd9384: begin digit0<=FOUR; digit1<=EIGHT; digit2<=THREE; digit3<=NINE; end
      16'd9385: begin digit0<=FIVE; digit1<=EIGHT; digit2<=THREE; digit3<=NINE; end
      16'd9386: begin digit0<=SIX; digit1<=EIGHT; digit2<=THREE; digit3<=NINE; end
      16'd9387: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=THREE; digit3<=NINE; end
      16'd9388: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=THREE; digit3<=NINE; end
      16'd9389: begin digit0<=NINE; digit1<=EIGHT; digit2<=THREE; digit3<=NINE; end
      16'd9390: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=NINE; end
      16'd9391: begin digit0<=ONE; digit1<=NINE; digit2<=THREE; digit3<=NINE; end
      16'd9392: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=NINE; end
      16'd9393: begin digit0<=THREE; digit1<=NINE; digit2<=THREE; digit3<=NINE; end
      16'd9394: begin digit0<=FOUR; digit1<=NINE; digit2<=THREE; digit3<=NINE; end
      16'd9395: begin digit0<=FIVE; digit1<=NINE; digit2<=THREE; digit3<=NINE; end
      16'd9396: begin digit0<=SIX; digit1<=NINE; digit2<=THREE; digit3<=NINE; end
      16'd9397: begin digit0<=SEVEN; digit1<=NINE; digit2<=THREE; digit3<=NINE; end
      16'd9398: begin digit0<=EIGHT; digit1<=NINE; digit2<=THREE; digit3<=NINE; end
      16'd9399: begin digit0<=NINE; digit1<=NINE; digit2<=THREE; digit3<=NINE; end
	  16'd9400: begin digit0<=ZERO; digit1<=ZERO; digit2<=FOUR; digit3<=NINE; end
      16'd9401: begin digit0<=ONE; digit1<=ZERO; digit2<=FOUR; digit3<=NINE; end
      16'd9402: begin digit0<=TWO; digit1<=ZERO; digit2<=FOUR; digit3<=NINE; end
      16'd9403: begin digit0<=THREE; digit1<=ZERO; digit2<=FOUR; digit3<=NINE; end
      16'd9404: begin digit0<=FOUR; digit1<=ZERO; digit2<=FOUR; digit3<=NINE; end
      16'd9405: begin digit0<=FIVE; digit1<=ZERO; digit2<=FOUR; digit3<=NINE; end
      16'd9406: begin digit0<=SIX; digit1<=ZERO; digit2<=FOUR; digit3<=NINE; end
      16'd9407: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FOUR; digit3<=NINE; end
      16'd9408: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FOUR; digit3<=NINE; end
      16'd9409: begin digit0<=NINE; digit1<=ZERO; digit2<=FOUR; digit3<=NINE; end
      16'd9410: begin digit0<=ZERO; digit1<=ONE; digit2<=FOUR; digit3<=NINE; end
      16'd9411: begin digit0<=ONE; digit1<=ONE; digit2<=FOUR; digit3<=NINE; end
      16'd9412: begin digit0<=TWO; digit1<=ONE; digit2<=FOUR; digit3<=NINE; end
      16'd9413: begin digit0<=THREE; digit1<=ONE; digit2<=FOUR; digit3<=NINE; end
      16'd9414: begin digit0<=FOUR; digit1<=ONE; digit2<=FOUR; digit3<=NINE; end
      16'd9415: begin digit0<=FIVE; digit1<=ONE; digit2<=FOUR; digit3<=NINE; end
      16'd9416: begin digit0<=SIX; digit1<=ONE; digit2<=FOUR; digit3<=NINE; end
      16'd9417: begin digit0<=SEVEN; digit1<=ONE; digit2<=FOUR; digit3<=NINE; end
      16'd9418: begin digit0<=EIGHT; digit1<=ONE; digit2<=FOUR; digit3<=NINE; end
      16'd9419: begin digit0<=NINE; digit1<=ONE; digit2<=FOUR; digit3<=NINE; end
      16'd9420: begin digit0<=ZERO; digit1<=TWO; digit2<=FOUR; digit3<=NINE; end
      16'd9421: begin digit0<=ONE; digit1<=TWO; digit2<=FOUR; digit3<=NINE; end
      16'd9422: begin digit0<=TWO; digit1<=TWO; digit2<=FOUR; digit3<=NINE; end
      16'd9423: begin digit0<=THREE; digit1<=TWO; digit2<=FOUR; digit3<=NINE; end
      16'd9424: begin digit0<=FOUR; digit1<=TWO; digit2<=FOUR; digit3<=NINE; end
      16'd9425: begin digit0<=FIVE; digit1<=TWO; digit2<=FOUR; digit3<=NINE; end
      16'd9426: begin digit0<=SIX; digit1<=TWO; digit2<=FOUR; digit3<=NINE; end
      16'd9427: begin digit0<=SEVEN; digit1<=TWO; digit2<=FOUR; digit3<=NINE; end
      16'd9428: begin digit0<=EIGHT; digit1<=TWO; digit2<=FOUR; digit3<=NINE; end
      16'd9429: begin digit0<=NINE; digit1<=TWO; digit2<=FOUR; digit3<=NINE; end
      16'd9430: begin digit0<=ZERO; digit1<=THREE; digit2<=FOUR; digit3<=NINE; end
      16'd9431: begin digit0<=ONE; digit1<=THREE; digit2<=FOUR; digit3<=NINE; end
      16'd9432: begin digit0<=TWO; digit1<=THREE; digit2<=FOUR; digit3<=NINE; end
      16'd9433: begin digit0<=THREE; digit1<=THREE; digit2<=FOUR; digit3<=NINE; end
      16'd9434: begin digit0<=FOUR; digit1<=THREE; digit2<=FOUR; digit3<=NINE; end
      16'd9435: begin digit0<=FIVE; digit1<=THREE; digit2<=FOUR; digit3<=NINE; end
      16'd9436: begin digit0<=SIX; digit1<=THREE; digit2<=FOUR; digit3<=NINE; end
      16'd9437: begin digit0<=SEVEN; digit1<=THREE; digit2<=FOUR; digit3<=NINE; end
      16'd9438: begin digit0<=EIGHT; digit1<=THREE; digit2<=FOUR; digit3<=NINE; end
      16'd9439: begin digit0<=NINE; digit1<=THREE; digit2<=FOUR; digit3<=NINE; end
      16'd9440: begin digit0<=ZERO; digit1<=FOUR; digit2<=FOUR; digit3<=NINE; end
      16'd9441: begin digit0<=ONE; digit1<=FOUR; digit2<=FOUR; digit3<=NINE; end
      16'd9442: begin digit0<=TWO; digit1<=FOUR; digit2<=FOUR; digit3<=NINE; end
      16'd9443: begin digit0<=THREE; digit1<=FOUR; digit2<=FOUR; digit3<=NINE; end
      16'd9444: begin digit0<=FOUR; digit1<=FOUR; digit2<=FOUR; digit3<=NINE; end
      16'd9445: begin digit0<=FIVE; digit1<=FOUR; digit2<=FOUR; digit3<=NINE; end
      16'd9446: begin digit0<=SIX; digit1<=FOUR; digit2<=FOUR; digit3<=NINE; end
      16'd9447: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FOUR; digit3<=NINE; end
      16'd9448: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FOUR; digit3<=NINE; end
      16'd9449: begin digit0<=NINE; digit1<=FOUR; digit2<=FOUR; digit3<=NINE; end
      16'd9450: begin digit0<=ZERO; digit1<=FIVE; digit2<=FOUR; digit3<=NINE; end
      16'd9451: begin digit0<=ONE; digit1<=FIVE; digit2<=FOUR; digit3<=NINE; end
      16'd9452: begin digit0<=TWO; digit1<=FIVE; digit2<=FOUR; digit3<=NINE; end
      16'd9453: begin digit0<=THREE; digit1<=FIVE; digit2<=FOUR; digit3<=NINE; end
      16'd9454: begin digit0<=FOUR; digit1<=FIVE; digit2<=FOUR; digit3<=NINE; end
      16'd9455: begin digit0<=FIVE; digit1<=FIVE; digit2<=FOUR; digit3<=NINE; end
      16'd9456: begin digit0<=SIX; digit1<=FIVE; digit2<=FOUR; digit3<=NINE; end
      16'd9457: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FOUR; digit3<=NINE; end
      16'd9458: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FOUR; digit3<=NINE; end
      16'd9459: begin digit0<=NINE; digit1<=FIVE; digit2<=FOUR; digit3<=NINE; end
      16'd9460: begin digit0<=ZERO; digit1<=SIX; digit2<=FOUR; digit3<=NINE; end
      16'd9461: begin digit0<=ONE; digit1<=SIX; digit2<=FOUR; digit3<=NINE; end
      16'd9462: begin digit0<=TWO; digit1<=SIX; digit2<=FOUR; digit3<=NINE; end
      16'd9463: begin digit0<=THREE; digit1<=SIX; digit2<=FOUR; digit3<=NINE; end
      16'd9464: begin digit0<=FOUR; digit1<=SIX; digit2<=FOUR; digit3<=NINE; end
      16'd9465: begin digit0<=FIVE; digit1<=SIX; digit2<=FOUR; digit3<=NINE; end
      16'd9466: begin digit0<=SIX; digit1<=SIX; digit2<=FOUR; digit3<=NINE; end
      16'd9467: begin digit0<=SEVEN; digit1<=SIX; digit2<=FOUR; digit3<=NINE; end
      16'd9468: begin digit0<=EIGHT; digit1<=SIX; digit2<=FOUR; digit3<=NINE; end
      16'd9469: begin digit0<=NINE; digit1<=SIX; digit2<=FOUR; digit3<=NINE; end
      16'd9470: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FOUR; digit3<=NINE; end
      16'd9471: begin digit0<=ONE; digit1<=SEVEN; digit2<=FOUR; digit3<=NINE; end
      16'd9472: begin digit0<=TWO; digit1<=SEVEN; digit2<=FOUR; digit3<=NINE; end
      16'd9473: begin digit0<=THREE; digit1<=SEVEN; digit2<=FOUR; digit3<=NINE; end
      16'd9474: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FOUR; digit3<=NINE; end
      16'd9475: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FOUR; digit3<=NINE; end
      16'd9476: begin digit0<=SIX; digit1<=SEVEN; digit2<=FOUR; digit3<=NINE; end
      16'd9477: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FOUR; digit3<=NINE; end
      16'd9478: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FOUR; digit3<=NINE; end
      16'd9479: begin digit0<=NINE; digit1<=SEVEN; digit2<=FOUR; digit3<=NINE; end
      16'd9480: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=NINE; end
      16'd9481: begin digit0<=ONE; digit1<=EIGHT; digit2<=FOUR; digit3<=NINE; end
      16'd9482: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=NINE; end
      16'd9483: begin digit0<=THREE; digit1<=EIGHT; digit2<=FOUR; digit3<=NINE; end
      16'd9484: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FOUR; digit3<=NINE; end
      16'd9485: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FOUR; digit3<=NINE; end
      16'd9486: begin digit0<=SIX; digit1<=EIGHT; digit2<=FOUR; digit3<=NINE; end
      16'd9487: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FOUR; digit3<=NINE; end
      16'd9488: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FOUR; digit3<=NINE; end
      16'd9489: begin digit0<=NINE; digit1<=EIGHT; digit2<=FOUR; digit3<=NINE; end
      16'd9490: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=NINE; end
      16'd9491: begin digit0<=ONE; digit1<=NINE; digit2<=FOUR; digit3<=NINE; end
      16'd9492: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=NINE; end
      16'd9493: begin digit0<=THREE; digit1<=NINE; digit2<=FOUR; digit3<=NINE; end
      16'd9494: begin digit0<=FOUR; digit1<=NINE; digit2<=FOUR; digit3<=NINE; end
      16'd9495: begin digit0<=FIVE; digit1<=NINE; digit2<=FOUR; digit3<=NINE; end
      16'd9496: begin digit0<=SIX; digit1<=NINE; digit2<=FOUR; digit3<=NINE; end
      16'd9497: begin digit0<=SEVEN; digit1<=NINE; digit2<=FOUR; digit3<=NINE; end
      16'd9498: begin digit0<=EIGHT; digit1<=NINE; digit2<=FOUR; digit3<=NINE; end
      16'd9499: begin digit0<=NINE; digit1<=NINE; digit2<=FOUR; digit3<=NINE; end
	  16'd9500: begin digit0<=ZERO; digit1<=ZERO; digit2<=FIVE; digit3<=NINE; end
      16'd9501: begin digit0<=ONE; digit1<=ZERO; digit2<=FIVE; digit3<=NINE; end
      16'd9502: begin digit0<=TWO; digit1<=ZERO; digit2<=FIVE; digit3<=NINE; end
      16'd9503: begin digit0<=THREE; digit1<=ZERO; digit2<=FIVE; digit3<=NINE; end
      16'd9504: begin digit0<=FOUR; digit1<=ZERO; digit2<=FIVE; digit3<=NINE; end
      16'd9505: begin digit0<=FIVE; digit1<=ZERO; digit2<=FIVE; digit3<=NINE; end
      16'd9506: begin digit0<=SIX; digit1<=ZERO; digit2<=FIVE; digit3<=NINE; end
      16'd9507: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FIVE; digit3<=NINE; end
      16'd9508: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FIVE; digit3<=NINE; end
      16'd9509: begin digit0<=NINE; digit1<=ZERO; digit2<=FIVE; digit3<=NINE; end
      16'd9510: begin digit0<=ZERO; digit1<=ONE; digit2<=FIVE; digit3<=NINE; end
      16'd9511: begin digit0<=ONE; digit1<=ONE; digit2<=FIVE; digit3<=NINE; end
      16'd9512: begin digit0<=TWO; digit1<=ONE; digit2<=FIVE; digit3<=NINE; end
      16'd9513: begin digit0<=THREE; digit1<=ONE; digit2<=FIVE; digit3<=NINE; end
      16'd9514: begin digit0<=FOUR; digit1<=ONE; digit2<=FIVE; digit3<=NINE; end
      16'd9515: begin digit0<=FIVE; digit1<=ONE; digit2<=FIVE; digit3<=NINE; end
      16'd9516: begin digit0<=SIX; digit1<=ONE; digit2<=FIVE; digit3<=NINE; end
      16'd9517: begin digit0<=SEVEN; digit1<=ONE; digit2<=FIVE; digit3<=NINE; end
      16'd9518: begin digit0<=EIGHT; digit1<=ONE; digit2<=FIVE; digit3<=NINE; end
      16'd9519: begin digit0<=NINE; digit1<=ONE; digit2<=FIVE; digit3<=NINE; end
      16'd9520: begin digit0<=ZERO; digit1<=TWO; digit2<=FIVE; digit3<=NINE; end
      16'd9521: begin digit0<=ONE; digit1<=TWO; digit2<=FIVE; digit3<=NINE; end
      16'd9522: begin digit0<=TWO; digit1<=TWO; digit2<=FIVE; digit3<=NINE; end
      16'd9523: begin digit0<=THREE; digit1<=TWO; digit2<=FIVE; digit3<=NINE; end
      16'd9524: begin digit0<=FOUR; digit1<=TWO; digit2<=FIVE; digit3<=NINE; end
      16'd9525: begin digit0<=FIVE; digit1<=TWO; digit2<=FIVE; digit3<=NINE; end
      16'd9526: begin digit0<=SIX; digit1<=TWO; digit2<=FIVE; digit3<=NINE; end
      16'd9527: begin digit0<=SEVEN; digit1<=TWO; digit2<=FIVE; digit3<=NINE; end
      16'd9528: begin digit0<=EIGHT; digit1<=TWO; digit2<=FIVE; digit3<=NINE; end
      16'd9529: begin digit0<=NINE; digit1<=TWO; digit2<=FIVE; digit3<=NINE; end
      16'd9530: begin digit0<=ZERO; digit1<=THREE; digit2<=FIVE; digit3<=NINE; end
      16'd9531: begin digit0<=ONE; digit1<=THREE; digit2<=FIVE; digit3<=NINE; end
      16'd9532: begin digit0<=TWO; digit1<=THREE; digit2<=FIVE; digit3<=NINE; end
      16'd9533: begin digit0<=THREE; digit1<=THREE; digit2<=FIVE; digit3<=NINE; end
      16'd9534: begin digit0<=FOUR; digit1<=THREE; digit2<=FIVE; digit3<=NINE; end
      16'd9535: begin digit0<=FIVE; digit1<=THREE; digit2<=FIVE; digit3<=NINE; end
      16'd9536: begin digit0<=SIX; digit1<=THREE; digit2<=FIVE; digit3<=NINE; end
      16'd9537: begin digit0<=SEVEN; digit1<=THREE; digit2<=FIVE; digit3<=NINE; end
      16'd9538: begin digit0<=EIGHT; digit1<=THREE; digit2<=FIVE; digit3<=NINE; end
      16'd9539: begin digit0<=NINE; digit1<=THREE; digit2<=FIVE; digit3<=NINE; end
      16'd9540: begin digit0<=ZERO; digit1<=FOUR; digit2<=FIVE; digit3<=NINE; end
      16'd9541: begin digit0<=ONE; digit1<=FOUR; digit2<=FIVE; digit3<=NINE; end
      16'd9542: begin digit0<=TWO; digit1<=FOUR; digit2<=FIVE; digit3<=NINE; end
      16'd9543: begin digit0<=THREE; digit1<=FOUR; digit2<=FIVE; digit3<=NINE; end
      16'd9544: begin digit0<=FOUR; digit1<=FOUR; digit2<=FIVE; digit3<=NINE; end
      16'd9545: begin digit0<=FIVE; digit1<=FOUR; digit2<=FIVE; digit3<=NINE; end
      16'd9546: begin digit0<=SIX; digit1<=FOUR; digit2<=FIVE; digit3<=NINE; end
      16'd9547: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FIVE; digit3<=NINE; end
      16'd9548: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FIVE; digit3<=NINE; end
      16'd9549: begin digit0<=NINE; digit1<=FOUR; digit2<=FIVE; digit3<=NINE; end
      16'd9550: begin digit0<=ZERO; digit1<=FIVE; digit2<=FIVE; digit3<=NINE; end
      16'd9551: begin digit0<=ONE; digit1<=FIVE; digit2<=FIVE; digit3<=NINE; end
      16'd9552: begin digit0<=TWO; digit1<=FIVE; digit2<=FIVE; digit3<=NINE; end
      16'd9553: begin digit0<=THREE; digit1<=FIVE; digit2<=FIVE; digit3<=NINE; end
      16'd9554: begin digit0<=FOUR; digit1<=FIVE; digit2<=FIVE; digit3<=NINE; end
      16'd9555: begin digit0<=FIVE; digit1<=FIVE; digit2<=FIVE; digit3<=NINE; end
      16'd9556: begin digit0<=SIX; digit1<=FIVE; digit2<=FIVE; digit3<=NINE; end
      16'd9557: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FIVE; digit3<=NINE; end
      16'd9558: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FIVE; digit3<=NINE; end
      16'd9559: begin digit0<=NINE; digit1<=FIVE; digit2<=FIVE; digit3<=NINE; end
      16'd9560: begin digit0<=ZERO; digit1<=SIX; digit2<=FIVE; digit3<=NINE; end
      16'd9561: begin digit0<=ONE; digit1<=SIX; digit2<=FIVE; digit3<=NINE; end
      16'd9562: begin digit0<=TWO; digit1<=SIX; digit2<=FIVE; digit3<=NINE; end
      16'd9563: begin digit0<=THREE; digit1<=SIX; digit2<=FIVE; digit3<=NINE; end
      16'd9564: begin digit0<=FOUR; digit1<=SIX; digit2<=FIVE; digit3<=NINE; end
      16'd9565: begin digit0<=FIVE; digit1<=SIX; digit2<=FIVE; digit3<=NINE; end
      16'd9566: begin digit0<=SIX; digit1<=SIX; digit2<=FIVE; digit3<=NINE; end
      16'd9567: begin digit0<=SEVEN; digit1<=SIX; digit2<=FIVE; digit3<=NINE; end
      16'd9568: begin digit0<=EIGHT; digit1<=SIX; digit2<=FIVE; digit3<=NINE; end
      16'd9569: begin digit0<=NINE; digit1<=SIX; digit2<=FIVE; digit3<=NINE; end
      16'd9570: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FIVE; digit3<=NINE; end
      16'd9571: begin digit0<=ONE; digit1<=SEVEN; digit2<=FIVE; digit3<=NINE; end
      16'd9572: begin digit0<=TWO; digit1<=SEVEN; digit2<=FIVE; digit3<=NINE; end
      16'd9573: begin digit0<=THREE; digit1<=SEVEN; digit2<=FIVE; digit3<=NINE; end
      16'd9574: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FIVE; digit3<=NINE; end
      16'd9575: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FIVE; digit3<=NINE; end
      16'd9576: begin digit0<=SIX; digit1<=SEVEN; digit2<=FIVE; digit3<=NINE; end
      16'd9577: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FIVE; digit3<=NINE; end
      16'd9578: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FIVE; digit3<=NINE; end
      16'd9579: begin digit0<=NINE; digit1<=SEVEN; digit2<=FIVE; digit3<=NINE; end
      16'd9580: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=NINE; end
      16'd9581: begin digit0<=ONE; digit1<=EIGHT; digit2<=FIVE; digit3<=NINE; end
      16'd9582: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=NINE; end
      16'd9583: begin digit0<=THREE; digit1<=EIGHT; digit2<=FIVE; digit3<=NINE; end
      16'd9584: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FIVE; digit3<=NINE; end
      16'd9585: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FIVE; digit3<=NINE; end
      16'd9586: begin digit0<=SIX; digit1<=EIGHT; digit2<=FIVE; digit3<=NINE; end
      16'd9587: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FIVE; digit3<=NINE; end
      16'd9588: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FIVE; digit3<=NINE; end
      16'd9589: begin digit0<=NINE; digit1<=EIGHT; digit2<=FIVE; digit3<=NINE; end
      16'd9590: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=NINE; end
      16'd9591: begin digit0<=ONE; digit1<=NINE; digit2<=FIVE; digit3<=NINE; end
      16'd9592: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=NINE; end
      16'd9593: begin digit0<=THREE; digit1<=NINE; digit2<=FIVE; digit3<=NINE; end
      16'd9594: begin digit0<=FOUR; digit1<=NINE; digit2<=FIVE; digit3<=NINE; end
      16'd9595: begin digit0<=FIVE; digit1<=NINE; digit2<=FIVE; digit3<=NINE; end
      16'd9596: begin digit0<=SIX; digit1<=NINE; digit2<=FIVE; digit3<=NINE; end
      16'd9597: begin digit0<=SEVEN; digit1<=NINE; digit2<=FIVE; digit3<=NINE; end
      16'd9598: begin digit0<=EIGHT; digit1<=NINE; digit2<=FIVE; digit3<=NINE; end
      16'd9599: begin digit0<=NINE; digit1<=NINE; digit2<=FIVE; digit3<=NINE; end
	  16'd9600: begin digit0<=ZERO; digit1<=ZERO; digit2<=SIX; digit3<=NINE; end
      16'd9601: begin digit0<=ONE; digit1<=ZERO; digit2<=SIX; digit3<=NINE; end
      16'd9602: begin digit0<=TWO; digit1<=ZERO; digit2<=SIX; digit3<=NINE; end
      16'd9603: begin digit0<=THREE; digit1<=ZERO; digit2<=SIX; digit3<=NINE; end
      16'd9604: begin digit0<=FOUR; digit1<=ZERO; digit2<=SIX; digit3<=NINE; end
      16'd9605: begin digit0<=FIVE; digit1<=ZERO; digit2<=SIX; digit3<=NINE; end
      16'd9606: begin digit0<=SIX; digit1<=ZERO; digit2<=SIX; digit3<=NINE; end
      16'd9607: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SIX; digit3<=NINE; end
      16'd9608: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SIX; digit3<=NINE; end
      16'd9609: begin digit0<=NINE; digit1<=ZERO; digit2<=SIX; digit3<=NINE; end
      16'd9610: begin digit0<=ZERO; digit1<=ONE; digit2<=SIX; digit3<=NINE; end
      16'd9611: begin digit0<=ONE; digit1<=ONE; digit2<=SIX; digit3<=NINE; end
      16'd9612: begin digit0<=TWO; digit1<=ONE; digit2<=SIX; digit3<=NINE; end
      16'd9613: begin digit0<=THREE; digit1<=ONE; digit2<=SIX; digit3<=NINE; end
      16'd9614: begin digit0<=FOUR; digit1<=ONE; digit2<=SIX; digit3<=NINE; end
      16'd9615: begin digit0<=FIVE; digit1<=ONE; digit2<=SIX; digit3<=NINE; end
      16'd9616: begin digit0<=SIX; digit1<=ONE; digit2<=SIX; digit3<=NINE; end
      16'd9617: begin digit0<=SEVEN; digit1<=ONE; digit2<=SIX; digit3<=NINE; end
      16'd9618: begin digit0<=EIGHT; digit1<=ONE; digit2<=SIX; digit3<=NINE; end
      16'd9619: begin digit0<=NINE; digit1<=ONE; digit2<=SIX; digit3<=NINE; end
      16'd9620: begin digit0<=ZERO; digit1<=TWO; digit2<=SIX; digit3<=NINE; end
      16'd9621: begin digit0<=ONE; digit1<=TWO; digit2<=SIX; digit3<=NINE; end
      16'd9622: begin digit0<=TWO; digit1<=TWO; digit2<=SIX; digit3<=NINE; end
      16'd9623: begin digit0<=THREE; digit1<=TWO; digit2<=SIX; digit3<=NINE; end
      16'd9624: begin digit0<=FOUR; digit1<=TWO; digit2<=SIX; digit3<=NINE; end
      16'd9625: begin digit0<=FIVE; digit1<=TWO; digit2<=SIX; digit3<=NINE; end
      16'd9626: begin digit0<=SIX; digit1<=TWO; digit2<=SIX; digit3<=NINE; end
      16'd9627: begin digit0<=SEVEN; digit1<=TWO; digit2<=SIX; digit3<=NINE; end
      16'd9628: begin digit0<=EIGHT; digit1<=TWO; digit2<=SIX; digit3<=NINE; end
      16'd9629: begin digit0<=NINE; digit1<=TWO; digit2<=SIX; digit3<=NINE; end
      16'd9630: begin digit0<=ZERO; digit1<=THREE; digit2<=SIX; digit3<=NINE; end
      16'd9631: begin digit0<=ONE; digit1<=THREE; digit2<=SIX; digit3<=NINE; end
      16'd9632: begin digit0<=TWO; digit1<=THREE; digit2<=SIX; digit3<=NINE; end
      16'd9633: begin digit0<=THREE; digit1<=THREE; digit2<=SIX; digit3<=NINE; end
      16'd9634: begin digit0<=FOUR; digit1<=THREE; digit2<=SIX; digit3<=NINE; end
      16'd9635: begin digit0<=FIVE; digit1<=THREE; digit2<=SIX; digit3<=NINE; end
      16'd9636: begin digit0<=SIX; digit1<=THREE; digit2<=SIX; digit3<=NINE; end
      16'd9637: begin digit0<=SEVEN; digit1<=THREE; digit2<=SIX; digit3<=NINE; end
      16'd9638: begin digit0<=EIGHT; digit1<=THREE; digit2<=SIX; digit3<=NINE; end
      16'd9639: begin digit0<=NINE; digit1<=THREE; digit2<=SIX; digit3<=NINE; end
      16'd9640: begin digit0<=ZERO; digit1<=FOUR; digit2<=SIX; digit3<=NINE; end
      16'd9641: begin digit0<=ONE; digit1<=FOUR; digit2<=SIX; digit3<=NINE; end
      16'd9642: begin digit0<=TWO; digit1<=FOUR; digit2<=SIX; digit3<=NINE; end
      16'd9643: begin digit0<=THREE; digit1<=FOUR; digit2<=SIX; digit3<=NINE; end
      16'd9644: begin digit0<=FOUR; digit1<=FOUR; digit2<=SIX; digit3<=NINE; end
      16'd9645: begin digit0<=FIVE; digit1<=FOUR; digit2<=SIX; digit3<=NINE; end
      16'd9646: begin digit0<=SIX; digit1<=FOUR; digit2<=SIX; digit3<=NINE; end
      16'd9647: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SIX; digit3<=NINE; end
      16'd9648: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SIX; digit3<=NINE; end
      16'd9649: begin digit0<=NINE; digit1<=FOUR; digit2<=SIX; digit3<=NINE; end
      16'd9650: begin digit0<=ZERO; digit1<=FIVE; digit2<=SIX; digit3<=NINE; end
      16'd9651: begin digit0<=ONE; digit1<=FIVE; digit2<=SIX; digit3<=NINE; end
      16'd9652: begin digit0<=TWO; digit1<=FIVE; digit2<=SIX; digit3<=NINE; end
      16'd9653: begin digit0<=THREE; digit1<=FIVE; digit2<=SIX; digit3<=NINE; end
      16'd9654: begin digit0<=FOUR; digit1<=FIVE; digit2<=SIX; digit3<=NINE; end
      16'd9655: begin digit0<=FIVE; digit1<=FIVE; digit2<=SIX; digit3<=NINE; end
      16'd9656: begin digit0<=SIX; digit1<=FIVE; digit2<=SIX; digit3<=NINE; end
      16'd9657: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SIX; digit3<=NINE; end
      16'd9658: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SIX; digit3<=NINE; end
      16'd9659: begin digit0<=NINE; digit1<=FIVE; digit2<=SIX; digit3<=NINE; end
      16'd9660: begin digit0<=ZERO; digit1<=SIX; digit2<=SIX; digit3<=NINE; end
      16'd9661: begin digit0<=ONE; digit1<=SIX; digit2<=SIX; digit3<=NINE; end
      16'd9662: begin digit0<=TWO; digit1<=SIX; digit2<=SIX; digit3<=NINE; end
      16'd9663: begin digit0<=THREE; digit1<=SIX; digit2<=SIX; digit3<=NINE; end
      16'd9664: begin digit0<=FOUR; digit1<=SIX; digit2<=SIX; digit3<=NINE; end
      16'd9665: begin digit0<=FIVE; digit1<=SIX; digit2<=SIX; digit3<=NINE; end
      16'd9666: begin digit0<=SIX; digit1<=SIX; digit2<=SIX; digit3<=NINE; end
      16'd9667: begin digit0<=SEVEN; digit1<=SIX; digit2<=SIX; digit3<=NINE; end
      16'd9668: begin digit0<=EIGHT; digit1<=SIX; digit2<=SIX; digit3<=NINE; end
      16'd9669: begin digit0<=NINE; digit1<=SIX; digit2<=SIX; digit3<=NINE; end
      16'd9670: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SIX; digit3<=NINE; end
      16'd9671: begin digit0<=ONE; digit1<=SEVEN; digit2<=SIX; digit3<=NINE; end
      16'd9672: begin digit0<=TWO; digit1<=SEVEN; digit2<=SIX; digit3<=NINE; end
      16'd9673: begin digit0<=THREE; digit1<=SEVEN; digit2<=SIX; digit3<=NINE; end
      16'd9674: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SIX; digit3<=NINE; end
      16'd9675: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SIX; digit3<=NINE; end
      16'd9676: begin digit0<=SIX; digit1<=SEVEN; digit2<=SIX; digit3<=NINE; end
      16'd9677: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SIX; digit3<=NINE; end
      16'd9678: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SIX; digit3<=NINE; end
      16'd9679: begin digit0<=NINE; digit1<=SEVEN; digit2<=SIX; digit3<=NINE; end
      16'd9680: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=NINE; end
      16'd9681: begin digit0<=ONE; digit1<=EIGHT; digit2<=SIX; digit3<=NINE; end
      16'd9682: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=NINE; end
      16'd9683: begin digit0<=THREE; digit1<=EIGHT; digit2<=SIX; digit3<=NINE; end
      16'd9684: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SIX; digit3<=NINE; end
      16'd9685: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SIX; digit3<=NINE; end
      16'd9686: begin digit0<=SIX; digit1<=EIGHT; digit2<=SIX; digit3<=NINE; end
      16'd9687: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SIX; digit3<=NINE; end
      16'd9688: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SIX; digit3<=NINE; end
      16'd9689: begin digit0<=NINE; digit1<=EIGHT; digit2<=SIX; digit3<=NINE; end
      16'd9690: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=NINE; end
      16'd9691: begin digit0<=ONE; digit1<=NINE; digit2<=SIX; digit3<=NINE; end
      16'd9692: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=NINE; end
      16'd9693: begin digit0<=THREE; digit1<=NINE; digit2<=SIX; digit3<=NINE; end
      16'd9694: begin digit0<=FOUR; digit1<=NINE; digit2<=SIX; digit3<=NINE; end
      16'd9695: begin digit0<=FIVE; digit1<=NINE; digit2<=SIX; digit3<=NINE; end
      16'd9696: begin digit0<=SIX; digit1<=NINE; digit2<=SIX; digit3<=NINE; end
      16'd9697: begin digit0<=SEVEN; digit1<=NINE; digit2<=SIX; digit3<=NINE; end
      16'd9698: begin digit0<=EIGHT; digit1<=NINE; digit2<=SIX; digit3<=NINE; end
      16'd9699: begin digit0<=NINE; digit1<=NINE; digit2<=SIX; digit3<=NINE; end
	  16'd9700: begin digit0<=ZERO; digit1<=ZERO; digit2<=SEVEN; digit3<=NINE; end
      16'd9701: begin digit0<=ONE; digit1<=ZERO; digit2<=SEVEN; digit3<=NINE; end
      16'd9702: begin digit0<=TWO; digit1<=ZERO; digit2<=SEVEN; digit3<=NINE; end
      16'd9703: begin digit0<=THREE; digit1<=ZERO; digit2<=SEVEN; digit3<=NINE; end
      16'd9704: begin digit0<=FOUR; digit1<=ZERO; digit2<=SEVEN; digit3<=NINE; end
      16'd9705: begin digit0<=FIVE; digit1<=ZERO; digit2<=SEVEN; digit3<=NINE; end
      16'd9706: begin digit0<=SIX; digit1<=ZERO; digit2<=SEVEN; digit3<=NINE; end
      16'd9707: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SEVEN; digit3<=NINE; end
      16'd9708: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SEVEN; digit3<=NINE; end
      16'd9709: begin digit0<=NINE; digit1<=ZERO; digit2<=SEVEN; digit3<=NINE; end
      16'd9710: begin digit0<=ZERO; digit1<=ONE; digit2<=SEVEN; digit3<=NINE; end
      16'd9711: begin digit0<=ONE; digit1<=ONE; digit2<=SEVEN; digit3<=NINE; end
      16'd9712: begin digit0<=TWO; digit1<=ONE; digit2<=SEVEN; digit3<=NINE; end
      16'd9713: begin digit0<=THREE; digit1<=ONE; digit2<=SEVEN; digit3<=NINE; end
      16'd9714: begin digit0<=FOUR; digit1<=ONE; digit2<=SEVEN; digit3<=NINE; end
      16'd9715: begin digit0<=FIVE; digit1<=ONE; digit2<=SEVEN; digit3<=NINE; end
      16'd9716: begin digit0<=SIX; digit1<=ONE; digit2<=SEVEN; digit3<=NINE; end
      16'd9717: begin digit0<=SEVEN; digit1<=ONE; digit2<=SEVEN; digit3<=NINE; end
      16'd9718: begin digit0<=EIGHT; digit1<=ONE; digit2<=SEVEN; digit3<=NINE; end
      16'd9719: begin digit0<=NINE; digit1<=ONE; digit2<=SEVEN; digit3<=NINE; end
      16'd9720: begin digit0<=ZERO; digit1<=TWO; digit2<=SEVEN; digit3<=NINE; end
      16'd9721: begin digit0<=ONE; digit1<=TWO; digit2<=SEVEN; digit3<=NINE; end
      16'd9722: begin digit0<=TWO; digit1<=TWO; digit2<=SEVEN; digit3<=NINE; end
      16'd9723: begin digit0<=THREE; digit1<=TWO; digit2<=SEVEN; digit3<=NINE; end
      16'd9724: begin digit0<=FOUR; digit1<=TWO; digit2<=SEVEN; digit3<=NINE; end
      16'd9725: begin digit0<=FIVE; digit1<=TWO; digit2<=SEVEN; digit3<=NINE; end
      16'd9726: begin digit0<=SIX; digit1<=TWO; digit2<=SEVEN; digit3<=NINE; end
      16'd9727: begin digit0<=SEVEN; digit1<=TWO; digit2<=SEVEN; digit3<=NINE; end
      16'd9728: begin digit0<=EIGHT; digit1<=TWO; digit2<=SEVEN; digit3<=NINE; end
      16'd9729: begin digit0<=NINE; digit1<=TWO; digit2<=SEVEN; digit3<=NINE; end
      16'd9730: begin digit0<=ZERO; digit1<=THREE; digit2<=SEVEN; digit3<=NINE; end
      16'd9731: begin digit0<=ONE; digit1<=THREE; digit2<=SEVEN; digit3<=NINE; end
      16'd9732: begin digit0<=TWO; digit1<=THREE; digit2<=SEVEN; digit3<=NINE; end
      16'd9733: begin digit0<=THREE; digit1<=THREE; digit2<=SEVEN; digit3<=NINE; end
      16'd9734: begin digit0<=FOUR; digit1<=THREE; digit2<=SEVEN; digit3<=NINE; end
      16'd9735: begin digit0<=FIVE; digit1<=THREE; digit2<=SEVEN; digit3<=NINE; end
      16'd9736: begin digit0<=SIX; digit1<=THREE; digit2<=SEVEN; digit3<=NINE; end
      16'd9737: begin digit0<=SEVEN; digit1<=THREE; digit2<=SEVEN; digit3<=NINE; end
      16'd9738: begin digit0<=EIGHT; digit1<=THREE; digit2<=SEVEN; digit3<=NINE; end
      16'd9739: begin digit0<=NINE; digit1<=THREE; digit2<=SEVEN; digit3<=NINE; end
      16'd9740: begin digit0<=ZERO; digit1<=FOUR; digit2<=SEVEN; digit3<=NINE; end
      16'd9741: begin digit0<=ONE; digit1<=FOUR; digit2<=SEVEN; digit3<=NINE; end
      16'd9742: begin digit0<=TWO; digit1<=FOUR; digit2<=SEVEN; digit3<=NINE; end
      16'd9743: begin digit0<=THREE; digit1<=FOUR; digit2<=SEVEN; digit3<=NINE; end
      16'd9744: begin digit0<=FOUR; digit1<=FOUR; digit2<=SEVEN; digit3<=NINE; end
      16'd9745: begin digit0<=FIVE; digit1<=FOUR; digit2<=SEVEN; digit3<=NINE; end
      16'd9746: begin digit0<=SIX; digit1<=FOUR; digit2<=SEVEN; digit3<=NINE; end
      16'd9747: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SEVEN; digit3<=NINE; end
      16'd9748: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SEVEN; digit3<=NINE; end
      16'd9749: begin digit0<=NINE; digit1<=FOUR; digit2<=SEVEN; digit3<=NINE; end
      16'd9750: begin digit0<=ZERO; digit1<=FIVE; digit2<=SEVEN; digit3<=NINE; end
      16'd9751: begin digit0<=ONE; digit1<=FIVE; digit2<=SEVEN; digit3<=NINE; end
      16'd9752: begin digit0<=TWO; digit1<=FIVE; digit2<=SEVEN; digit3<=NINE; end
      16'd9753: begin digit0<=THREE; digit1<=FIVE; digit2<=SEVEN; digit3<=NINE; end
      16'd9754: begin digit0<=FOUR; digit1<=FIVE; digit2<=SEVEN; digit3<=NINE; end
      16'd9755: begin digit0<=FIVE; digit1<=FIVE; digit2<=SEVEN; digit3<=NINE; end
      16'd9756: begin digit0<=SIX; digit1<=FIVE; digit2<=SEVEN; digit3<=NINE; end
      16'd9757: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SEVEN; digit3<=NINE; end
      16'd9758: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SEVEN; digit3<=NINE; end
      16'd9759: begin digit0<=NINE; digit1<=FIVE; digit2<=SEVEN; digit3<=NINE; end
      16'd9760: begin digit0<=ZERO; digit1<=SIX; digit2<=SEVEN; digit3<=NINE; end
      16'd9761: begin digit0<=ONE; digit1<=SIX; digit2<=SEVEN; digit3<=NINE; end
      16'd9762: begin digit0<=TWO; digit1<=SIX; digit2<=SEVEN; digit3<=NINE; end
      16'd9763: begin digit0<=THREE; digit1<=SIX; digit2<=SEVEN; digit3<=NINE; end
      16'd9764: begin digit0<=FOUR; digit1<=SIX; digit2<=SEVEN; digit3<=NINE; end
      16'd9765: begin digit0<=FIVE; digit1<=SIX; digit2<=SEVEN; digit3<=NINE; end
      16'd9766: begin digit0<=SIX; digit1<=SIX; digit2<=SEVEN; digit3<=NINE; end
      16'd9767: begin digit0<=SEVEN; digit1<=SIX; digit2<=SEVEN; digit3<=NINE; end
      16'd9768: begin digit0<=EIGHT; digit1<=SIX; digit2<=SEVEN; digit3<=NINE; end
      16'd9769: begin digit0<=NINE; digit1<=SIX; digit2<=SEVEN; digit3<=NINE; end
      16'd9770: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SEVEN; digit3<=NINE; end
      16'd9771: begin digit0<=ONE; digit1<=SEVEN; digit2<=SEVEN; digit3<=NINE; end
      16'd9772: begin digit0<=TWO; digit1<=SEVEN; digit2<=SEVEN; digit3<=NINE; end
      16'd9773: begin digit0<=THREE; digit1<=SEVEN; digit2<=SEVEN; digit3<=NINE; end
      16'd9774: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SEVEN; digit3<=NINE; end
      16'd9775: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SEVEN; digit3<=NINE; end
      16'd9776: begin digit0<=SIX; digit1<=SEVEN; digit2<=SEVEN; digit3<=NINE; end
      16'd9777: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SEVEN; digit3<=NINE; end
      16'd9778: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SEVEN; digit3<=NINE; end
      16'd9779: begin digit0<=NINE; digit1<=SEVEN; digit2<=SEVEN; digit3<=NINE; end
      16'd9780: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=NINE; end
      16'd9781: begin digit0<=ONE; digit1<=EIGHT; digit2<=SEVEN; digit3<=NINE; end
      16'd9782: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=NINE; end
      16'd9783: begin digit0<=THREE; digit1<=EIGHT; digit2<=SEVEN; digit3<=NINE; end
      16'd9784: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SEVEN; digit3<=NINE; end
      16'd9785: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SEVEN; digit3<=NINE; end
      16'd9786: begin digit0<=SIX; digit1<=EIGHT; digit2<=SEVEN; digit3<=NINE; end
      16'd9787: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SEVEN; digit3<=NINE; end
      16'd9788: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SEVEN; digit3<=NINE; end
      16'd9789: begin digit0<=NINE; digit1<=EIGHT; digit2<=SEVEN; digit3<=NINE; end
      16'd9790: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=NINE; end
      16'd9791: begin digit0<=ONE; digit1<=NINE; digit2<=SEVEN; digit3<=NINE; end
      16'd9792: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=NINE; end
      16'd9793: begin digit0<=THREE; digit1<=NINE; digit2<=SEVEN; digit3<=NINE; end
      16'd9794: begin digit0<=FOUR; digit1<=NINE; digit2<=SEVEN; digit3<=NINE; end
      16'd9795: begin digit0<=FIVE; digit1<=NINE; digit2<=SEVEN; digit3<=NINE; end
      16'd9796: begin digit0<=SIX; digit1<=NINE; digit2<=SEVEN; digit3<=NINE; end
      16'd9797: begin digit0<=SEVEN; digit1<=NINE; digit2<=SEVEN; digit3<=NINE; end
      16'd9798: begin digit0<=EIGHT; digit1<=NINE; digit2<=SEVEN; digit3<=NINE; end
      16'd9799: begin digit0<=NINE; digit1<=NINE; digit2<=SEVEN; digit3<=NINE; end
	  16'd9800: begin digit0<=ZERO; digit1<=ZERO; digit2<=EIGHT; digit3<=NINE; end
      16'd9801: begin digit0<=ONE; digit1<=ZERO; digit2<=EIGHT; digit3<=NINE; end
      16'd9802: begin digit0<=TWO; digit1<=ZERO; digit2<=EIGHT; digit3<=NINE; end
      16'd9803: begin digit0<=THREE; digit1<=ZERO; digit2<=EIGHT; digit3<=NINE; end
      16'd9804: begin digit0<=FOUR; digit1<=ZERO; digit2<=EIGHT; digit3<=NINE; end
      16'd9805: begin digit0<=FIVE; digit1<=ZERO; digit2<=EIGHT; digit3<=NINE; end
      16'd9806: begin digit0<=SIX; digit1<=ZERO; digit2<=EIGHT; digit3<=NINE; end
      16'd9807: begin digit0<=SEVEN; digit1<=ZERO; digit2<=EIGHT; digit3<=NINE; end
      16'd9808: begin digit0<=EIGHT; digit1<=ZERO; digit2<=EIGHT; digit3<=NINE; end
      16'd9809: begin digit0<=NINE; digit1<=ZERO; digit2<=EIGHT; digit3<=NINE; end
      16'd9810: begin digit0<=ZERO; digit1<=ONE; digit2<=EIGHT; digit3<=NINE; end
      16'd9811: begin digit0<=ONE; digit1<=ONE; digit2<=EIGHT; digit3<=NINE; end
      16'd9812: begin digit0<=TWO; digit1<=ONE; digit2<=EIGHT; digit3<=NINE; end
      16'd9813: begin digit0<=THREE; digit1<=ONE; digit2<=EIGHT; digit3<=NINE; end
      16'd9814: begin digit0<=FOUR; digit1<=ONE; digit2<=EIGHT; digit3<=NINE; end
      16'd9815: begin digit0<=FIVE; digit1<=ONE; digit2<=EIGHT; digit3<=NINE; end
      16'd9816: begin digit0<=SIX; digit1<=ONE; digit2<=EIGHT; digit3<=NINE; end
      16'd9817: begin digit0<=SEVEN; digit1<=ONE; digit2<=EIGHT; digit3<=NINE; end
      16'd9818: begin digit0<=EIGHT; digit1<=ONE; digit2<=EIGHT; digit3<=NINE; end
      16'd9819: begin digit0<=NINE; digit1<=ONE; digit2<=EIGHT; digit3<=NINE; end
      16'd9820: begin digit0<=ZERO; digit1<=TWO; digit2<=EIGHT; digit3<=NINE; end
      16'd9821: begin digit0<=ONE; digit1<=TWO; digit2<=EIGHT; digit3<=NINE; end
      16'd9822: begin digit0<=TWO; digit1<=TWO; digit2<=EIGHT; digit3<=NINE; end
      16'd9823: begin digit0<=THREE; digit1<=TWO; digit2<=EIGHT; digit3<=NINE; end
      16'd9824: begin digit0<=FOUR; digit1<=TWO; digit2<=EIGHT; digit3<=NINE; end
      16'd9825: begin digit0<=FIVE; digit1<=TWO; digit2<=EIGHT; digit3<=NINE; end
      16'd9826: begin digit0<=SIX; digit1<=TWO; digit2<=EIGHT; digit3<=NINE; end
      16'd9827: begin digit0<=SEVEN; digit1<=TWO; digit2<=EIGHT; digit3<=NINE; end
      16'd9828: begin digit0<=EIGHT; digit1<=TWO; digit2<=EIGHT; digit3<=NINE; end
      16'd9829: begin digit0<=NINE; digit1<=TWO; digit2<=EIGHT; digit3<=NINE; end
      16'd9830: begin digit0<=ZERO; digit1<=THREE; digit2<=EIGHT; digit3<=NINE; end
      16'd9831: begin digit0<=ONE; digit1<=THREE; digit2<=EIGHT; digit3<=NINE; end
      16'd9832: begin digit0<=TWO; digit1<=THREE; digit2<=EIGHT; digit3<=NINE; end
      16'd9833: begin digit0<=THREE; digit1<=THREE; digit2<=EIGHT; digit3<=NINE; end
      16'd9834: begin digit0<=FOUR; digit1<=THREE; digit2<=EIGHT; digit3<=NINE; end
      16'd9835: begin digit0<=FIVE; digit1<=THREE; digit2<=EIGHT; digit3<=NINE; end
      16'd9836: begin digit0<=SIX; digit1<=THREE; digit2<=EIGHT; digit3<=NINE; end
      16'd9837: begin digit0<=SEVEN; digit1<=THREE; digit2<=EIGHT; digit3<=NINE; end
      16'd9838: begin digit0<=EIGHT; digit1<=THREE; digit2<=EIGHT; digit3<=NINE; end
      16'd9839: begin digit0<=NINE; digit1<=THREE; digit2<=EIGHT; digit3<=NINE; end
      16'd9840: begin digit0<=ZERO; digit1<=FOUR; digit2<=EIGHT; digit3<=NINE; end
      16'd9841: begin digit0<=ONE; digit1<=FOUR; digit2<=EIGHT; digit3<=NINE; end
      16'd9842: begin digit0<=TWO; digit1<=FOUR; digit2<=EIGHT; digit3<=NINE; end
      16'd9843: begin digit0<=THREE; digit1<=FOUR; digit2<=EIGHT; digit3<=NINE; end
      16'd9844: begin digit0<=FOUR; digit1<=FOUR; digit2<=EIGHT; digit3<=NINE; end
      16'd9845: begin digit0<=FIVE; digit1<=FOUR; digit2<=EIGHT; digit3<=NINE; end
      16'd9846: begin digit0<=SIX; digit1<=FOUR; digit2<=EIGHT; digit3<=NINE; end
      16'd9847: begin digit0<=SEVEN; digit1<=FOUR; digit2<=EIGHT; digit3<=NINE; end
      16'd9848: begin digit0<=EIGHT; digit1<=FOUR; digit2<=EIGHT; digit3<=NINE; end
      16'd9849: begin digit0<=NINE; digit1<=FOUR; digit2<=EIGHT; digit3<=NINE; end
      16'd9850: begin digit0<=ZERO; digit1<=FIVE; digit2<=EIGHT; digit3<=NINE; end
      16'd9851: begin digit0<=ONE; digit1<=FIVE; digit2<=EIGHT; digit3<=NINE; end
      16'd9852: begin digit0<=TWO; digit1<=FIVE; digit2<=EIGHT; digit3<=NINE; end
      16'd9853: begin digit0<=THREE; digit1<=FIVE; digit2<=EIGHT; digit3<=NINE; end
      16'd9854: begin digit0<=FOUR; digit1<=FIVE; digit2<=EIGHT; digit3<=NINE; end
      16'd9855: begin digit0<=FIVE; digit1<=FIVE; digit2<=EIGHT; digit3<=NINE; end
      16'd9856: begin digit0<=SIX; digit1<=FIVE; digit2<=EIGHT; digit3<=NINE; end
      16'd9857: begin digit0<=SEVEN; digit1<=FIVE; digit2<=EIGHT; digit3<=NINE; end
      16'd9858: begin digit0<=EIGHT; digit1<=FIVE; digit2<=EIGHT; digit3<=NINE; end
      16'd9859: begin digit0<=NINE; digit1<=FIVE; digit2<=EIGHT; digit3<=NINE; end
      16'd9860: begin digit0<=ZERO; digit1<=SIX; digit2<=EIGHT; digit3<=NINE; end
      16'd9861: begin digit0<=ONE; digit1<=SIX; digit2<=EIGHT; digit3<=NINE; end
      16'd9862: begin digit0<=TWO; digit1<=SIX; digit2<=EIGHT; digit3<=NINE; end
      16'd9863: begin digit0<=THREE; digit1<=SIX; digit2<=EIGHT; digit3<=NINE; end
      16'd9864: begin digit0<=FOUR; digit1<=SIX; digit2<=EIGHT; digit3<=NINE; end
      16'd9865: begin digit0<=FIVE; digit1<=SIX; digit2<=EIGHT; digit3<=NINE; end
      16'd9866: begin digit0<=SIX; digit1<=SIX; digit2<=EIGHT; digit3<=NINE; end
      16'd9867: begin digit0<=SEVEN; digit1<=SIX; digit2<=EIGHT; digit3<=NINE; end
      16'd9868: begin digit0<=EIGHT; digit1<=SIX; digit2<=EIGHT; digit3<=NINE; end
      16'd9869: begin digit0<=NINE; digit1<=SIX; digit2<=EIGHT; digit3<=NINE; end
      16'd9870: begin digit0<=ZERO; digit1<=SEVEN; digit2<=EIGHT; digit3<=NINE; end
      16'd9871: begin digit0<=ONE; digit1<=SEVEN; digit2<=EIGHT; digit3<=NINE; end
      16'd9872: begin digit0<=TWO; digit1<=SEVEN; digit2<=EIGHT; digit3<=NINE; end
      16'd9873: begin digit0<=THREE; digit1<=SEVEN; digit2<=EIGHT; digit3<=NINE; end
      16'd9874: begin digit0<=FOUR; digit1<=SEVEN; digit2<=EIGHT; digit3<=NINE; end
      16'd9875: begin digit0<=FIVE; digit1<=SEVEN; digit2<=EIGHT; digit3<=NINE; end
      16'd9876: begin digit0<=SIX; digit1<=SEVEN; digit2<=EIGHT; digit3<=NINE; end
      16'd9877: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=EIGHT; digit3<=NINE; end
      16'd9878: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=EIGHT; digit3<=NINE; end
      16'd9879: begin digit0<=NINE; digit1<=SEVEN; digit2<=EIGHT; digit3<=NINE; end
      16'd9880: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=NINE; end
      16'd9881: begin digit0<=ONE; digit1<=EIGHT; digit2<=EIGHT; digit3<=NINE; end
      16'd9882: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=NINE; end
      16'd9883: begin digit0<=THREE; digit1<=EIGHT; digit2<=EIGHT; digit3<=NINE; end
      16'd9884: begin digit0<=FOUR; digit1<=EIGHT; digit2<=EIGHT; digit3<=NINE; end
      16'd9885: begin digit0<=FIVE; digit1<=EIGHT; digit2<=EIGHT; digit3<=NINE; end
      16'd9886: begin digit0<=SIX; digit1<=EIGHT; digit2<=EIGHT; digit3<=NINE; end
      16'd9887: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=EIGHT; digit3<=NINE; end
      16'd9888: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=EIGHT; digit3<=NINE; end
      16'd9889: begin digit0<=NINE; digit1<=EIGHT; digit2<=EIGHT; digit3<=NINE; end
      16'd9890: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=NINE; end
      16'd9891: begin digit0<=ONE; digit1<=NINE; digit2<=EIGHT; digit3<=NINE; end
      16'd9892: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=NINE; end
      16'd9893: begin digit0<=THREE; digit1<=NINE; digit2<=EIGHT; digit3<=NINE; end
      16'd9894: begin digit0<=FOUR; digit1<=NINE; digit2<=EIGHT; digit3<=NINE; end
      16'd9895: begin digit0<=FIVE; digit1<=NINE; digit2<=EIGHT; digit3<=NINE; end
      16'd9896: begin digit0<=SIX; digit1<=NINE; digit2<=EIGHT; digit3<=NINE; end
      16'd9897: begin digit0<=SEVEN; digit1<=NINE; digit2<=EIGHT; digit3<=NINE; end
      16'd9898: begin digit0<=EIGHT; digit1<=NINE; digit2<=EIGHT; digit3<=NINE; end
      16'd9899: begin digit0<=NINE; digit1<=NINE; digit2<=EIGHT; digit3<=NINE; end
	  16'd9900: begin digit0<=ZERO; digit1<=ZERO; digit2<=NINE; digit3<=NINE; end
      16'd9901: begin digit0<=ONE; digit1<=ZERO; digit2<=NINE; digit3<=NINE; end
      16'd9902: begin digit0<=TWO; digit1<=ZERO; digit2<=NINE; digit3<=NINE; end
      16'd9903: begin digit0<=THREE; digit1<=ZERO; digit2<=NINE; digit3<=NINE; end
      16'd9904: begin digit0<=FOUR; digit1<=ZERO; digit2<=NINE; digit3<=NINE; end
      16'd9905: begin digit0<=FIVE; digit1<=ZERO; digit2<=NINE; digit3<=NINE; end
      16'd9906: begin digit0<=SIX; digit1<=ZERO; digit2<=NINE; digit3<=NINE; end
      16'd9907: begin digit0<=SEVEN; digit1<=ZERO; digit2<=NINE; digit3<=NINE; end
      16'd9908: begin digit0<=EIGHT; digit1<=ZERO; digit2<=NINE; digit3<=NINE; end
      16'd9909: begin digit0<=NINE; digit1<=ZERO; digit2<=NINE; digit3<=NINE; end
      16'd9910: begin digit0<=ZERO; digit1<=ONE; digit2<=NINE; digit3<=NINE; end
      16'd9911: begin digit0<=ONE; digit1<=ONE; digit2<=NINE; digit3<=NINE; end
      16'd9912: begin digit0<=TWO; digit1<=ONE; digit2<=NINE; digit3<=NINE; end
      16'd9913: begin digit0<=THREE; digit1<=ONE; digit2<=NINE; digit3<=NINE; end
      16'd9914: begin digit0<=FOUR; digit1<=ONE; digit2<=NINE; digit3<=NINE; end
      16'd9915: begin digit0<=FIVE; digit1<=ONE; digit2<=NINE; digit3<=NINE; end
      16'd9916: begin digit0<=SIX; digit1<=ONE; digit2<=NINE; digit3<=NINE; end
      16'd9917: begin digit0<=SEVEN; digit1<=ONE; digit2<=NINE; digit3<=NINE; end
      16'd9918: begin digit0<=EIGHT; digit1<=ONE; digit2<=NINE; digit3<=NINE; end
      16'd9919: begin digit0<=NINE; digit1<=ONE; digit2<=NINE; digit3<=NINE; end
      16'd9920: begin digit0<=ZERO; digit1<=TWO; digit2<=NINE; digit3<=NINE; end
      16'd9921: begin digit0<=ONE; digit1<=TWO; digit2<=NINE; digit3<=NINE; end
      16'd9922: begin digit0<=TWO; digit1<=TWO; digit2<=NINE; digit3<=NINE; end
      16'd9923: begin digit0<=THREE; digit1<=TWO; digit2<=NINE; digit3<=NINE; end
      16'd9924: begin digit0<=FOUR; digit1<=TWO; digit2<=NINE; digit3<=NINE; end
      16'd9925: begin digit0<=FIVE; digit1<=TWO; digit2<=NINE; digit3<=NINE; end
      16'd9926: begin digit0<=SIX; digit1<=TWO; digit2<=NINE; digit3<=NINE; end
      16'd9927: begin digit0<=SEVEN; digit1<=TWO; digit2<=NINE; digit3<=NINE; end
      16'd9928: begin digit0<=EIGHT; digit1<=TWO; digit2<=NINE; digit3<=NINE; end
      16'd9929: begin digit0<=NINE; digit1<=TWO; digit2<=NINE; digit3<=NINE; end
      16'd9930: begin digit0<=ZERO; digit1<=THREE; digit2<=NINE; digit3<=NINE; end
      16'd9931: begin digit0<=ONE; digit1<=THREE; digit2<=NINE; digit3<=NINE; end
      16'd9932: begin digit0<=TWO; digit1<=THREE; digit2<=NINE; digit3<=NINE; end
      16'd9933: begin digit0<=THREE; digit1<=THREE; digit2<=NINE; digit3<=NINE; end
      16'd9934: begin digit0<=FOUR; digit1<=THREE; digit2<=NINE; digit3<=NINE; end
      16'd9935: begin digit0<=FIVE; digit1<=THREE; digit2<=NINE; digit3<=NINE; end
      16'd9936: begin digit0<=SIX; digit1<=THREE; digit2<=NINE; digit3<=NINE; end
      16'd9937: begin digit0<=SEVEN; digit1<=THREE; digit2<=NINE; digit3<=NINE; end
      16'd9938: begin digit0<=EIGHT; digit1<=THREE; digit2<=NINE; digit3<=NINE; end
      16'd9939: begin digit0<=NINE; digit1<=THREE; digit2<=NINE; digit3<=NINE; end
      16'd9940: begin digit0<=ZERO; digit1<=FOUR; digit2<=NINE; digit3<=NINE; end
      16'd9941: begin digit0<=ONE; digit1<=FOUR; digit2<=NINE; digit3<=NINE; end
      16'd9942: begin digit0<=TWO; digit1<=FOUR; digit2<=NINE; digit3<=NINE; end
      16'd9943: begin digit0<=THREE; digit1<=FOUR; digit2<=NINE; digit3<=NINE; end
      16'd9944: begin digit0<=FOUR; digit1<=FOUR; digit2<=NINE; digit3<=NINE; end
      16'd9945: begin digit0<=FIVE; digit1<=FOUR; digit2<=NINE; digit3<=NINE; end
      16'd9946: begin digit0<=SIX; digit1<=FOUR; digit2<=NINE; digit3<=NINE; end
      16'd9947: begin digit0<=SEVEN; digit1<=FOUR; digit2<=NINE; digit3<=NINE; end
      16'd9948: begin digit0<=EIGHT; digit1<=FOUR; digit2<=NINE; digit3<=NINE; end
      16'd9949: begin digit0<=NINE; digit1<=FOUR; digit2<=NINE; digit3<=NINE; end
      16'd9950: begin digit0<=ZERO; digit1<=FIVE; digit2<=NINE; digit3<=NINE; end
      16'd9951: begin digit0<=ONE; digit1<=FIVE; digit2<=NINE; digit3<=NINE; end
      16'd9952: begin digit0<=TWO; digit1<=FIVE; digit2<=NINE; digit3<=NINE; end
      16'd9953: begin digit0<=THREE; digit1<=FIVE; digit2<=NINE; digit3<=NINE; end
      16'd9954: begin digit0<=FOUR; digit1<=FIVE; digit2<=NINE; digit3<=NINE; end
      16'd9955: begin digit0<=FIVE; digit1<=FIVE; digit2<=NINE; digit3<=NINE; end
      16'd9956: begin digit0<=SIX; digit1<=FIVE; digit2<=NINE; digit3<=NINE; end
      16'd9957: begin digit0<=SEVEN; digit1<=FIVE; digit2<=NINE; digit3<=NINE; end
      16'd9958: begin digit0<=EIGHT; digit1<=FIVE; digit2<=NINE; digit3<=NINE; end
      16'd9959: begin digit0<=NINE; digit1<=FIVE; digit2<=NINE; digit3<=NINE; end
      16'd9960: begin digit0<=ZERO; digit1<=SIX; digit2<=NINE; digit3<=NINE; end
      16'd9961: begin digit0<=ONE; digit1<=SIX; digit2<=NINE; digit3<=NINE; end
      16'd9962: begin digit0<=TWO; digit1<=SIX; digit2<=NINE; digit3<=NINE; end
      16'd9963: begin digit0<=THREE; digit1<=SIX; digit2<=NINE; digit3<=NINE; end
      16'd9964: begin digit0<=FOUR; digit1<=SIX; digit2<=NINE; digit3<=NINE; end
      16'd9965: begin digit0<=FIVE; digit1<=SIX; digit2<=NINE; digit3<=NINE; end
      16'd9966: begin digit0<=SIX; digit1<=SIX; digit2<=NINE; digit3<=NINE; end
      16'd9967: begin digit0<=SEVEN; digit1<=SIX; digit2<=NINE; digit3<=NINE; end
      16'd9968: begin digit0<=EIGHT; digit1<=SIX; digit2<=NINE; digit3<=NINE; end
      16'd9969: begin digit0<=NINE; digit1<=SIX; digit2<=NINE; digit3<=NINE; end
      16'd9970: begin digit0<=ZERO; digit1<=SEVEN; digit2<=NINE; digit3<=NINE; end
      16'd9971: begin digit0<=ONE; digit1<=SEVEN; digit2<=NINE; digit3<=NINE; end
      16'd9972: begin digit0<=TWO; digit1<=SEVEN; digit2<=NINE; digit3<=NINE; end
      16'd9973: begin digit0<=THREE; digit1<=SEVEN; digit2<=NINE; digit3<=NINE; end
      16'd9974: begin digit0<=FOUR; digit1<=SEVEN; digit2<=NINE; digit3<=NINE; end
      16'd9975: begin digit0<=FIVE; digit1<=SEVEN; digit2<=NINE; digit3<=NINE; end
      16'd9976: begin digit0<=SIX; digit1<=SEVEN; digit2<=NINE; digit3<=NINE; end
      16'd9977: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=NINE; digit3<=NINE; end
      16'd9978: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=NINE; digit3<=NINE; end
      16'd9979: begin digit0<=NINE; digit1<=SEVEN; digit2<=NINE; digit3<=NINE; end
      16'd9980: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=NINE; end
      16'd9981: begin digit0<=ONE; digit1<=EIGHT; digit2<=NINE; digit3<=NINE; end
      16'd9982: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=NINE; end
      16'd9983: begin digit0<=THREE; digit1<=EIGHT; digit2<=NINE; digit3<=NINE; end
      16'd9984: begin digit0<=FOUR; digit1<=EIGHT; digit2<=NINE; digit3<=NINE; end
      16'd9985: begin digit0<=FIVE; digit1<=EIGHT; digit2<=NINE; digit3<=NINE; end
      16'd9986: begin digit0<=SIX; digit1<=EIGHT; digit2<=NINE; digit3<=NINE; end
      16'd9987: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=NINE; digit3<=NINE; end
      16'd9988: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=NINE; digit3<=NINE; end
      16'd9989: begin digit0<=NINE; digit1<=EIGHT; digit2<=NINE; digit3<=NINE; end
      16'd9990: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=NINE; end
      16'd9991: begin digit0<=ONE; digit1<=NINE; digit2<=NINE; digit3<=NINE; end
      16'd9992: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=NINE; end
      16'd9993: begin digit0<=THREE; digit1<=NINE; digit2<=NINE; digit3<=NINE; end
      16'd9994: begin digit0<=FOUR; digit1<=NINE; digit2<=NINE; digit3<=NINE; end
      16'd9995: begin digit0<=FIVE; digit1<=NINE; digit2<=NINE; digit3<=NINE; end
      16'd9996: begin digit0<=SIX; digit1<=NINE; digit2<=NINE; digit3<=NINE; end
      16'd9997: begin digit0<=SEVEN; digit1<=NINE; digit2<=NINE; digit3<=NINE; end
      16'd9998: begin digit0<=EIGHT; digit1<=NINE; digit2<=NINE; digit3<=NINE; end
      16'd9999: begin digit0<=NINE; digit1<=NINE; digit2<=NINE; digit3<=NINE; end
      default: begin digit0<=EMPTY; digit1<=EMPTY; digit2<=EMPTY; digit3<=EMPTY; end
    endcase
  else if (display_en & neg_en)
    case (tmp)
      16'd10000:begin digit0<=R; digit1<=R; digit2<=E; digit3<=EMPTY; end
      16'd0: begin digit0<=ZERO; digit1<=EMPTY; digit2<=EMPTY; digit3<=EMPTY; end
      16'd1: begin digit0<=ONE; digit1<=MIN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd2: begin digit0<=TWO; digit1<=MIN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd3: begin digit0<=THREE; digit1<=MIN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd4: begin digit0<=FOUR; digit1<=MIN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd5: begin digit0<=FIVE; digit1<=MIN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd6: begin digit0<=SIX; digit1<=MIN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd7: begin digit0<=SEVEN; digit1<=MIN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd8: begin digit0<=EIGHT; digit1<=MIN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd9: begin digit0<=NINE; digit1<=MIN; digit2<=EMPTY; digit3<=EMPTY; end
      16'd10: begin digit0<=ZERO; digit1<=ONE; digit2<=MIN; digit3<=EMPTY; end
      16'd11: begin digit0<=ONE; digit1<=ONE; digit2<=MIN; digit3<=EMPTY; end
      16'd12: begin digit0<=TWO; digit1<=ONE; digit2<=MIN; digit3<=EMPTY; end
      16'd13: begin digit0<=THREE; digit1<=ONE; digit2<=MIN; digit3<=EMPTY; end
      16'd14: begin digit0<=FOUR; digit1<=ONE; digit2<=MIN; digit3<=EMPTY; end
      16'd15: begin digit0<=FIVE; digit1<=ONE; digit2<=MIN; digit3<=EMPTY; end
      16'd16: begin digit0<=SIX; digit1<=ONE; digit2<=MIN; digit3<=EMPTY; end
      16'd17: begin digit0<=SEVEN; digit1<=ONE; digit2<=MIN; digit3<=EMPTY; end
      16'd18: begin digit0<=EIGHT; digit1<=ONE; digit2<=MIN; digit3<=EMPTY; end
      16'd19: begin digit0<=NINE; digit1<=ONE; digit2<=MIN; digit3<=EMPTY; end
      16'd20: begin digit0<=ZERO; digit1<=TWO; digit2<=MIN; digit3<=EMPTY; end
      16'd21: begin digit0<=ONE; digit1<=TWO; digit2<=MIN; digit3<=EMPTY; end
      16'd22: begin digit0<=TWO; digit1<=TWO; digit2<=MIN; digit3<=EMPTY; end
      16'd23: begin digit0<=THREE; digit1<=TWO; digit2<=MIN; digit3<=EMPTY; end
      16'd24: begin digit0<=FOUR; digit1<=TWO; digit2<=MIN; digit3<=EMPTY; end
      16'd25: begin digit0<=FIVE; digit1<=TWO; digit2<=MIN; digit3<=EMPTY; end
      16'd26: begin digit0<=SIX; digit1<=TWO; digit2<=MIN; digit3<=EMPTY; end
      16'd27: begin digit0<=SEVEN; digit1<=TWO; digit2<=MIN; digit3<=EMPTY; end
      16'd28: begin digit0<=EIGHT; digit1<=TWO; digit2<=MIN; digit3<=EMPTY; end
      16'd29: begin digit0<=NINE; digit1<=TWO; digit2<=MIN; digit3<=EMPTY; end
      16'd30: begin digit0<=ZERO; digit1<=THREE; digit2<=MIN; digit3<=EMPTY; end
      16'd31: begin digit0<=ONE; digit1<=THREE; digit2<=MIN; digit3<=EMPTY; end
      16'd32: begin digit0<=TWO; digit1<=THREE; digit2<=MIN; digit3<=EMPTY; end
      16'd33: begin digit0<=THREE; digit1<=THREE; digit2<=MIN; digit3<=EMPTY; end
      16'd34: begin digit0<=FOUR; digit1<=THREE; digit2<=MIN; digit3<=EMPTY; end
      16'd35: begin digit0<=FIVE; digit1<=THREE; digit2<=MIN; digit3<=EMPTY; end
      16'd36: begin digit0<=SIX; digit1<=THREE; digit2<=MIN; digit3<=EMPTY; end
      16'd37: begin digit0<=SEVEN; digit1<=THREE; digit2<=MIN; digit3<=EMPTY; end
      16'd38: begin digit0<=EIGHT; digit1<=THREE; digit2<=MIN; digit3<=EMPTY; end
      16'd39: begin digit0<=NINE; digit1<=THREE; digit2<=MIN; digit3<=EMPTY; end
      16'd40: begin digit0<=ZERO; digit1<=FOUR; digit2<=MIN; digit3<=EMPTY; end
      16'd41: begin digit0<=ONE; digit1<=FOUR; digit2<=MIN; digit3<=EMPTY; end
      16'd42: begin digit0<=TWO; digit1<=FOUR; digit2<=MIN; digit3<=EMPTY; end
      16'd43: begin digit0<=THREE; digit1<=FOUR; digit2<=MIN; digit3<=EMPTY; end
      16'd44: begin digit0<=FOUR; digit1<=FOUR; digit2<=MIN; digit3<=EMPTY; end
      16'd45: begin digit0<=FIVE; digit1<=FOUR; digit2<=MIN; digit3<=EMPTY; end
      16'd46: begin digit0<=SIX; digit1<=FOUR; digit2<=MIN; digit3<=EMPTY; end
      16'd47: begin digit0<=SEVEN; digit1<=FOUR; digit2<=MIN; digit3<=EMPTY; end
      16'd48: begin digit0<=EIGHT; digit1<=FOUR; digit2<=MIN; digit3<=EMPTY; end
      16'd49: begin digit0<=NINE; digit1<=FOUR; digit2<=MIN; digit3<=EMPTY; end
      16'd50: begin digit0<=ZERO; digit1<=FIVE; digit2<=MIN; digit3<=EMPTY; end
      16'd51: begin digit0<=ONE; digit1<=FIVE; digit2<=MIN; digit3<=EMPTY; end
      16'd52: begin digit0<=TWO; digit1<=FIVE; digit2<=MIN; digit3<=EMPTY; end
      16'd53: begin digit0<=THREE; digit1<=FIVE; digit2<=MIN; digit3<=EMPTY; end
      16'd54: begin digit0<=FOUR; digit1<=FIVE; digit2<=MIN; digit3<=EMPTY; end
      16'd55: begin digit0<=FIVE; digit1<=FIVE; digit2<=MIN; digit3<=EMPTY; end
      16'd56: begin digit0<=SIX; digit1<=FIVE; digit2<=MIN; digit3<=EMPTY; end
      16'd57: begin digit0<=SEVEN; digit1<=FIVE; digit2<=MIN; digit3<=EMPTY; end
      16'd58: begin digit0<=EIGHT; digit1<=FIVE; digit2<=MIN; digit3<=EMPTY; end
      16'd59: begin digit0<=NINE; digit1<=FIVE; digit2<=MIN; digit3<=EMPTY; end
      16'd60: begin digit0<=ZERO; digit1<=SIX; digit2<=MIN; digit3<=EMPTY; end
      16'd61: begin digit0<=ONE; digit1<=SIX; digit2<=MIN; digit3<=EMPTY; end
      16'd62: begin digit0<=TWO; digit1<=SIX; digit2<=MIN; digit3<=EMPTY; end
      16'd63: begin digit0<=THREE; digit1<=SIX; digit2<=MIN; digit3<=EMPTY; end
      16'd64: begin digit0<=FOUR; digit1<=SIX; digit2<=MIN; digit3<=EMPTY; end
      16'd65: begin digit0<=FIVE; digit1<=SIX; digit2<=MIN; digit3<=EMPTY; end
      16'd66: begin digit0<=SIX; digit1<=SIX; digit2<=MIN; digit3<=EMPTY; end
      16'd67: begin digit0<=SEVEN; digit1<=SIX; digit2<=MIN; digit3<=EMPTY; end
      16'd68: begin digit0<=EIGHT; digit1<=SIX; digit2<=MIN; digit3<=EMPTY; end
      16'd69: begin digit0<=NINE; digit1<=SIX; digit2<=MIN; digit3<=EMPTY; end
      16'd70: begin digit0<=ZERO; digit1<=SEVEN; digit2<=MIN; digit3<=EMPTY; end
      16'd71: begin digit0<=ONE; digit1<=SEVEN; digit2<=MIN; digit3<=EMPTY; end
      16'd72: begin digit0<=TWO; digit1<=SEVEN; digit2<=MIN; digit3<=EMPTY; end
      16'd73: begin digit0<=THREE; digit1<=SEVEN; digit2<=MIN; digit3<=EMPTY; end
      16'd74: begin digit0<=FOUR; digit1<=SEVEN; digit2<=MIN; digit3<=EMPTY; end
      16'd75: begin digit0<=FIVE; digit1<=SEVEN; digit2<=MIN; digit3<=EMPTY; end
      16'd76: begin digit0<=SIX; digit1<=SEVEN; digit2<=MIN; digit3<=EMPTY; end
      16'd77: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=MIN; digit3<=EMPTY; end
      16'd78: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=MIN; digit3<=EMPTY; end
      16'd79: begin digit0<=NINE; digit1<=SEVEN; digit2<=MIN; digit3<=EMPTY; end
      16'd80: begin digit0<=ZERO; digit1<=EIGHT; digit2<=MIN; digit3<=EMPTY; end
      16'd81: begin digit0<=ONE; digit1<=EIGHT; digit2<=MIN; digit3<=EMPTY; end
      16'd82: begin digit0<=ZERO; digit1<=EIGHT; digit2<=MIN; digit3<=EMPTY; end
      16'd83: begin digit0<=THREE; digit1<=EIGHT; digit2<=MIN; digit3<=EMPTY; end
      16'd84: begin digit0<=FOUR; digit1<=EIGHT; digit2<=MIN; digit3<=EMPTY; end
      16'd85: begin digit0<=FIVE; digit1<=EIGHT; digit2<=MIN; digit3<=EMPTY; end
      16'd86: begin digit0<=SIX; digit1<=EIGHT; digit2<=MIN; digit3<=EMPTY; end
      16'd87: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=MIN; digit3<=EMPTY; end
      16'd88: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=MIN; digit3<=EMPTY; end
      16'd89: begin digit0<=NINE; digit1<=EIGHT; digit2<=MIN; digit3<=EMPTY; end
      16'd90: begin digit0<=ZERO; digit1<=NINE; digit2<=MIN; digit3<=EMPTY; end
      16'd91: begin digit0<=ONE; digit1<=NINE; digit2<=MIN; digit3<=EMPTY; end
      16'd92: begin digit0<=ZERO; digit1<=NINE; digit2<=MIN; digit3<=EMPTY; end
      16'd93: begin digit0<=THREE; digit1<=NINE; digit2<=MIN; digit3<=EMPTY; end
      16'd94: begin digit0<=FOUR; digit1<=NINE; digit2<=MIN; digit3<=EMPTY; end
      16'd95: begin digit0<=FIVE; digit1<=NINE; digit2<=MIN; digit3<=EMPTY; end
      16'd96: begin digit0<=SIX; digit1<=NINE; digit2<=MIN; digit3<=EMPTY; end
      16'd97: begin digit0<=SEVEN; digit1<=NINE; digit2<=MIN; digit3<=EMPTY; end
      16'd98: begin digit0<=EIGHT; digit1<=NINE; digit2<=MIN; digit3<=EMPTY; end
      16'd99: begin digit0<=NINE; digit1<=NINE; digit2<=MIN; digit3<=EMPTY; end
	  16'd100: begin digit0<=ZERO; digit1<=ZERO; digit2<=ONE; digit3<=MIN; end
      16'd101: begin digit0<=ONE; digit1<=ZERO; digit2<=ONE; digit3<=MIN; end
      16'd102: begin digit0<=TWO; digit1<=ZERO; digit2<=ONE; digit3<=MIN; end
      16'd103: begin digit0<=THREE; digit1<=ZERO; digit2<=ONE; digit3<=MIN; end
      16'd104: begin digit0<=FOUR; digit1<=ZERO; digit2<=ONE; digit3<=MIN; end
      16'd105: begin digit0<=FIVE; digit1<=ZERO; digit2<=ONE; digit3<=MIN; end
      16'd106: begin digit0<=SIX; digit1<=ZERO; digit2<=ONE; digit3<=MIN; end
      16'd107: begin digit0<=SEVEN; digit1<=ZERO; digit2<=ONE; digit3<=MIN; end
      16'd108: begin digit0<=EIGHT; digit1<=ZERO; digit2<=ONE; digit3<=MIN; end
      16'd109: begin digit0<=NINE; digit1<=ZERO; digit2<=ONE; digit3<=MIN; end
      16'd110: begin digit0<=ZERO; digit1<=ONE; digit2<=ONE; digit3<=MIN; end
      16'd111: begin digit0<=ONE; digit1<=ONE; digit2<=ONE; digit3<=MIN; end
      16'd112: begin digit0<=TWO; digit1<=ONE; digit2<=ONE; digit3<=MIN; end
      16'd113: begin digit0<=THREE; digit1<=ONE; digit2<=ONE; digit3<=MIN; end
      16'd114: begin digit0<=FOUR; digit1<=ONE; digit2<=ONE; digit3<=MIN; end
      16'd115: begin digit0<=FIVE; digit1<=ONE; digit2<=ONE; digit3<=MIN; end
      16'd116: begin digit0<=SIX; digit1<=ONE; digit2<=ONE; digit3<=MIN; end
      16'd117: begin digit0<=SEVEN; digit1<=ONE; digit2<=ONE; digit3<=MIN; end
      16'd118: begin digit0<=EIGHT; digit1<=ONE; digit2<=ONE; digit3<=MIN; end
      16'd119: begin digit0<=NINE; digit1<=ONE; digit2<=ONE; digit3<=MIN; end
      16'd120: begin digit0<=ZERO; digit1<=TWO; digit2<=ONE; digit3<=MIN; end
      16'd121: begin digit0<=ONE; digit1<=TWO; digit2<=ONE; digit3<=MIN; end
      16'd122: begin digit0<=TWO; digit1<=TWO; digit2<=ONE; digit3<=MIN; end
      16'd123: begin digit0<=THREE; digit1<=TWO; digit2<=ONE; digit3<=MIN; end
      16'd124: begin digit0<=FOUR; digit1<=TWO; digit2<=ONE; digit3<=MIN; end
      16'd125: begin digit0<=FIVE; digit1<=TWO; digit2<=ONE; digit3<=MIN; end
      16'd126: begin digit0<=SIX; digit1<=TWO; digit2<=ONE; digit3<=MIN; end
      16'd127: begin digit0<=SEVEN; digit1<=TWO; digit2<=ONE; digit3<=MIN; end
      16'd128: begin digit0<=EIGHT; digit1<=TWO; digit2<=ONE; digit3<=MIN; end
      16'd129: begin digit0<=NINE; digit1<=TWO; digit2<=ONE; digit3<=MIN; end
      16'd130: begin digit0<=ZERO; digit1<=THREE; digit2<=ONE; digit3<=MIN; end
      16'd131: begin digit0<=ONE; digit1<=THREE; digit2<=ONE; digit3<=MIN; end
      16'd132: begin digit0<=TWO; digit1<=THREE; digit2<=ONE; digit3<=MIN; end
      16'd133: begin digit0<=THREE; digit1<=THREE; digit2<=ONE; digit3<=MIN; end
      16'd134: begin digit0<=FOUR; digit1<=THREE; digit2<=ONE; digit3<=MIN; end
      16'd135: begin digit0<=FIVE; digit1<=THREE; digit2<=ONE; digit3<=MIN; end
      16'd136: begin digit0<=SIX; digit1<=THREE; digit2<=ONE; digit3<=MIN; end
      16'd137: begin digit0<=SEVEN; digit1<=THREE; digit2<=ONE; digit3<=MIN; end
      16'd138: begin digit0<=EIGHT; digit1<=THREE; digit2<=ONE; digit3<=MIN; end
      16'd139: begin digit0<=NINE; digit1<=THREE; digit2<=ONE; digit3<=MIN; end
      16'd140: begin digit0<=ZERO; digit1<=FOUR; digit2<=ONE; digit3<=MIN; end
      16'd141: begin digit0<=ONE; digit1<=FOUR; digit2<=ONE; digit3<=MIN; end
      16'd142: begin digit0<=TWO; digit1<=FOUR; digit2<=ONE; digit3<=MIN; end
      16'd143: begin digit0<=THREE; digit1<=FOUR; digit2<=ONE; digit3<=MIN; end
      16'd144: begin digit0<=FOUR; digit1<=FOUR; digit2<=ONE; digit3<=MIN; end
      16'd145: begin digit0<=FIVE; digit1<=FOUR; digit2<=ONE; digit3<=MIN; end
      16'd146: begin digit0<=SIX; digit1<=FOUR; digit2<=ONE; digit3<=MIN; end
      16'd147: begin digit0<=SEVEN; digit1<=FOUR; digit2<=ONE; digit3<=MIN; end
      16'd148: begin digit0<=EIGHT; digit1<=FOUR; digit2<=ONE; digit3<=MIN; end
      16'd149: begin digit0<=NINE; digit1<=FOUR; digit2<=ONE; digit3<=MIN; end
      16'd150: begin digit0<=ZERO; digit1<=FIVE; digit2<=ONE; digit3<=MIN; end
      16'd151: begin digit0<=ONE; digit1<=FIVE; digit2<=ONE; digit3<=MIN; end
      16'd152: begin digit0<=TWO; digit1<=FIVE; digit2<=ONE; digit3<=MIN; end
      16'd153: begin digit0<=THREE; digit1<=FIVE; digit2<=ONE; digit3<=MIN; end
      16'd154: begin digit0<=FOUR; digit1<=FIVE; digit2<=ONE; digit3<=MIN; end
      16'd155: begin digit0<=FIVE; digit1<=FIVE; digit2<=ONE; digit3<=MIN; end
      16'd156: begin digit0<=SIX; digit1<=FIVE; digit2<=ONE; digit3<=MIN; end
      16'd157: begin digit0<=SEVEN; digit1<=FIVE; digit2<=ONE; digit3<=MIN; end
      16'd158: begin digit0<=EIGHT; digit1<=FIVE; digit2<=ONE; digit3<=MIN; end
      16'd159: begin digit0<=NINE; digit1<=FIVE; digit2<=ONE; digit3<=MIN; end
      16'd160: begin digit0<=ZERO; digit1<=SIX; digit2<=ONE; digit3<=MIN; end
      16'd161: begin digit0<=ONE; digit1<=SIX; digit2<=ONE; digit3<=MIN; end
      16'd162: begin digit0<=TWO; digit1<=SIX; digit2<=ONE; digit3<=MIN; end
      16'd163: begin digit0<=THREE; digit1<=SIX; digit2<=ONE; digit3<=MIN; end
      16'd164: begin digit0<=FOUR; digit1<=SIX; digit2<=ONE; digit3<=MIN; end
      16'd165: begin digit0<=FIVE; digit1<=SIX; digit2<=ONE; digit3<=MIN; end
      16'd166: begin digit0<=SIX; digit1<=SIX; digit2<=ONE; digit3<=MIN; end
      16'd167: begin digit0<=SEVEN; digit1<=SIX; digit2<=ONE; digit3<=MIN; end
      16'd168: begin digit0<=EIGHT; digit1<=SIX; digit2<=ONE; digit3<=MIN; end
      16'd169: begin digit0<=NINE; digit1<=SIX; digit2<=ONE; digit3<=MIN; end
      16'd170: begin digit0<=ZERO; digit1<=SEVEN; digit2<=ONE; digit3<=MIN; end
      16'd171: begin digit0<=ONE; digit1<=SEVEN; digit2<=ONE; digit3<=MIN; end
      16'd172: begin digit0<=TWO; digit1<=SEVEN; digit2<=ONE; digit3<=MIN; end
      16'd173: begin digit0<=THREE; digit1<=SEVEN; digit2<=ONE; digit3<=MIN; end
      16'd174: begin digit0<=FOUR; digit1<=SEVEN; digit2<=ONE; digit3<=MIN; end
      16'd175: begin digit0<=FIVE; digit1<=SEVEN; digit2<=ONE; digit3<=MIN; end
      16'd176: begin digit0<=SIX; digit1<=SEVEN; digit2<=ONE; digit3<=MIN; end
      16'd177: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=ONE; digit3<=MIN; end
      16'd178: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=ONE; digit3<=MIN; end
      16'd179: begin digit0<=NINE; digit1<=SEVEN; digit2<=ONE; digit3<=MIN; end
      16'd180: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=MIN; end
      16'd181: begin digit0<=ONE; digit1<=EIGHT; digit2<=ONE; digit3<=MIN; end
      16'd182: begin digit0<=ZERO; digit1<=EIGHT; digit2<=ONE; digit3<=MIN; end
      16'd183: begin digit0<=THREE; digit1<=EIGHT; digit2<=ONE; digit3<=MIN; end
      16'd184: begin digit0<=FOUR; digit1<=EIGHT; digit2<=ONE; digit3<=MIN; end
      16'd185: begin digit0<=FIVE; digit1<=EIGHT; digit2<=ONE; digit3<=MIN; end
      16'd186: begin digit0<=SIX; digit1<=EIGHT; digit2<=ONE; digit3<=MIN; end
      16'd187: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=ONE; digit3<=MIN; end
      16'd188: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=ONE; digit3<=MIN; end
      16'd189: begin digit0<=NINE; digit1<=EIGHT; digit2<=ONE; digit3<=MIN; end
      16'd190: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=MIN; end
      16'd191: begin digit0<=ONE; digit1<=NINE; digit2<=ONE; digit3<=MIN; end
      16'd192: begin digit0<=ZERO; digit1<=NINE; digit2<=ONE; digit3<=MIN; end
      16'd193: begin digit0<=THREE; digit1<=NINE; digit2<=ONE; digit3<=MIN; end
      16'd194: begin digit0<=FOUR; digit1<=NINE; digit2<=ONE; digit3<=MIN; end
      16'd195: begin digit0<=FIVE; digit1<=NINE; digit2<=ONE; digit3<=MIN; end
      16'd196: begin digit0<=SIX; digit1<=NINE; digit2<=ONE; digit3<=MIN; end
      16'd197: begin digit0<=SEVEN; digit1<=NINE; digit2<=ONE; digit3<=MIN; end
      16'd198: begin digit0<=EIGHT; digit1<=NINE; digit2<=ONE; digit3<=MIN; end
      16'd199: begin digit0<=NINE; digit1<=NINE; digit2<=ONE; digit3<=MIN; end
	  16'd200: begin digit0<=ZERO; digit1<=ZERO; digit2<=TWO; digit3<=MIN; end
      16'd201: begin digit0<=ONE; digit1<=ZERO; digit2<=TWO; digit3<=MIN; end
      16'd202: begin digit0<=TWO; digit1<=ZERO; digit2<=TWO; digit3<=MIN; end
      16'd203: begin digit0<=THREE; digit1<=ZERO; digit2<=TWO; digit3<=MIN; end
      16'd204: begin digit0<=FOUR; digit1<=ZERO; digit2<=TWO; digit3<=MIN; end
      16'd205: begin digit0<=FIVE; digit1<=ZERO; digit2<=TWO; digit3<=MIN; end
      16'd206: begin digit0<=SIX; digit1<=ZERO; digit2<=TWO; digit3<=MIN; end
      16'd207: begin digit0<=SEVEN; digit1<=ZERO; digit2<=TWO; digit3<=MIN; end
      16'd208: begin digit0<=EIGHT; digit1<=ZERO; digit2<=TWO; digit3<=MIN; end
      16'd209: begin digit0<=NINE; digit1<=ZERO; digit2<=TWO; digit3<=MIN; end
      16'd210: begin digit0<=ZERO; digit1<=ONE; digit2<=TWO; digit3<=MIN; end
      16'd211: begin digit0<=ONE; digit1<=ONE; digit2<=TWO; digit3<=MIN; end
      16'd212: begin digit0<=TWO; digit1<=ONE; digit2<=TWO; digit3<=MIN; end
      16'd213: begin digit0<=THREE; digit1<=ONE; digit2<=TWO; digit3<=MIN; end
      16'd214: begin digit0<=FOUR; digit1<=ONE; digit2<=TWO; digit3<=MIN; end
      16'd215: begin digit0<=FIVE; digit1<=ONE; digit2<=TWO; digit3<=MIN; end
      16'd216: begin digit0<=SIX; digit1<=ONE; digit2<=TWO; digit3<=MIN; end
      16'd217: begin digit0<=SEVEN; digit1<=ONE; digit2<=TWO; digit3<=MIN; end
      16'd218: begin digit0<=EIGHT; digit1<=ONE; digit2<=TWO; digit3<=MIN; end
      16'd219: begin digit0<=NINE; digit1<=ONE; digit2<=TWO; digit3<=MIN; end
      16'd220: begin digit0<=ZERO; digit1<=TWO; digit2<=TWO; digit3<=MIN; end
      16'd221: begin digit0<=ONE; digit1<=TWO; digit2<=TWO; digit3<=MIN; end
      16'd222: begin digit0<=TWO; digit1<=TWO; digit2<=TWO; digit3<=MIN; end
      16'd223: begin digit0<=THREE; digit1<=TWO; digit2<=TWO; digit3<=MIN; end
      16'd224: begin digit0<=FOUR; digit1<=TWO; digit2<=TWO; digit3<=MIN; end
      16'd225: begin digit0<=FIVE; digit1<=TWO; digit2<=TWO; digit3<=MIN; end
      16'd226: begin digit0<=SIX; digit1<=TWO; digit2<=TWO; digit3<=MIN; end
      16'd227: begin digit0<=SEVEN; digit1<=TWO; digit2<=TWO; digit3<=MIN; end
      16'd228: begin digit0<=EIGHT; digit1<=TWO; digit2<=TWO; digit3<=MIN; end
      16'd229: begin digit0<=NINE; digit1<=TWO; digit2<=TWO; digit3<=MIN; end
      16'd230: begin digit0<=ZERO; digit1<=THREE; digit2<=TWO; digit3<=MIN; end
      16'd231: begin digit0<=ONE; digit1<=THREE; digit2<=TWO; digit3<=MIN; end
      16'd232: begin digit0<=TWO; digit1<=THREE; digit2<=TWO; digit3<=MIN; end
      16'd233: begin digit0<=THREE; digit1<=THREE; digit2<=TWO; digit3<=MIN; end
      16'd234: begin digit0<=FOUR; digit1<=THREE; digit2<=TWO; digit3<=MIN; end
      16'd235: begin digit0<=FIVE; digit1<=THREE; digit2<=TWO; digit3<=MIN; end
      16'd236: begin digit0<=SIX; digit1<=THREE; digit2<=TWO; digit3<=MIN; end
      16'd237: begin digit0<=SEVEN; digit1<=THREE; digit2<=TWO; digit3<=MIN; end
      16'd238: begin digit0<=EIGHT; digit1<=THREE; digit2<=TWO; digit3<=MIN; end
      16'd239: begin digit0<=NINE; digit1<=THREE; digit2<=TWO; digit3<=MIN; end
      16'd240: begin digit0<=ZERO; digit1<=FOUR; digit2<=TWO; digit3<=MIN; end
      16'd241: begin digit0<=ONE; digit1<=FOUR; digit2<=TWO; digit3<=MIN; end
      16'd242: begin digit0<=TWO; digit1<=FOUR; digit2<=TWO; digit3<=MIN; end
      16'd243: begin digit0<=THREE; digit1<=FOUR; digit2<=TWO; digit3<=MIN; end
      16'd244: begin digit0<=FOUR; digit1<=FOUR; digit2<=TWO; digit3<=MIN; end
      16'd245: begin digit0<=FIVE; digit1<=FOUR; digit2<=TWO; digit3<=MIN; end
      16'd246: begin digit0<=SIX; digit1<=FOUR; digit2<=TWO; digit3<=MIN; end
      16'd247: begin digit0<=SEVEN; digit1<=FOUR; digit2<=TWO; digit3<=MIN; end
      16'd248: begin digit0<=EIGHT; digit1<=FOUR; digit2<=TWO; digit3<=MIN; end
      16'd249: begin digit0<=NINE; digit1<=FOUR; digit2<=TWO; digit3<=MIN; end
      16'd250: begin digit0<=ZERO; digit1<=FIVE; digit2<=TWO; digit3<=MIN; end
      16'd251: begin digit0<=ONE; digit1<=FIVE; digit2<=TWO; digit3<=MIN; end
      16'd252: begin digit0<=TWO; digit1<=FIVE; digit2<=TWO; digit3<=MIN; end
      16'd253: begin digit0<=THREE; digit1<=FIVE; digit2<=TWO; digit3<=MIN; end
      16'd254: begin digit0<=FOUR; digit1<=FIVE; digit2<=TWO; digit3<=MIN; end
      16'd255: begin digit0<=FIVE; digit1<=FIVE; digit2<=TWO; digit3<=MIN; end
      16'd256: begin digit0<=SIX; digit1<=FIVE; digit2<=TWO; digit3<=MIN; end
      16'd257: begin digit0<=SEVEN; digit1<=FIVE; digit2<=TWO; digit3<=MIN; end
      16'd258: begin digit0<=EIGHT; digit1<=FIVE; digit2<=TWO; digit3<=MIN; end
      16'd259: begin digit0<=NINE; digit1<=FIVE; digit2<=TWO; digit3<=MIN; end
      16'd260: begin digit0<=ZERO; digit1<=SIX; digit2<=TWO; digit3<=MIN; end
      16'd261: begin digit0<=ONE; digit1<=SIX; digit2<=TWO; digit3<=MIN; end
      16'd262: begin digit0<=TWO; digit1<=SIX; digit2<=TWO; digit3<=MIN; end
      16'd263: begin digit0<=THREE; digit1<=SIX; digit2<=TWO; digit3<=MIN; end
      16'd264: begin digit0<=FOUR; digit1<=SIX; digit2<=TWO; digit3<=MIN; end
      16'd265: begin digit0<=FIVE; digit1<=SIX; digit2<=TWO; digit3<=MIN; end
      16'd266: begin digit0<=SIX; digit1<=SIX; digit2<=TWO; digit3<=MIN; end
      16'd267: begin digit0<=SEVEN; digit1<=SIX; digit2<=TWO; digit3<=MIN; end
      16'd268: begin digit0<=EIGHT; digit1<=SIX; digit2<=TWO; digit3<=MIN; end
      16'd269: begin digit0<=NINE; digit1<=SIX; digit2<=TWO; digit3<=MIN; end
      16'd270: begin digit0<=ZERO; digit1<=SEVEN; digit2<=TWO; digit3<=MIN; end
      16'd271: begin digit0<=ONE; digit1<=SEVEN; digit2<=TWO; digit3<=MIN; end
      16'd272: begin digit0<=TWO; digit1<=SEVEN; digit2<=TWO; digit3<=MIN; end
      16'd273: begin digit0<=THREE; digit1<=SEVEN; digit2<=TWO; digit3<=MIN; end
      16'd274: begin digit0<=FOUR; digit1<=SEVEN; digit2<=TWO; digit3<=MIN; end
      16'd275: begin digit0<=FIVE; digit1<=SEVEN; digit2<=TWO; digit3<=MIN; end
      16'd276: begin digit0<=SIX; digit1<=SEVEN; digit2<=TWO; digit3<=MIN; end
      16'd277: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=TWO; digit3<=MIN; end
      16'd278: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=TWO; digit3<=MIN; end
      16'd279: begin digit0<=NINE; digit1<=SEVEN; digit2<=TWO; digit3<=MIN; end
      16'd280: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=MIN; end
      16'd281: begin digit0<=ONE; digit1<=EIGHT; digit2<=TWO; digit3<=MIN; end
      16'd282: begin digit0<=ZERO; digit1<=EIGHT; digit2<=TWO; digit3<=MIN; end
      16'd283: begin digit0<=THREE; digit1<=EIGHT; digit2<=TWO; digit3<=MIN; end
      16'd284: begin digit0<=FOUR; digit1<=EIGHT; digit2<=TWO; digit3<=MIN; end
      16'd285: begin digit0<=FIVE; digit1<=EIGHT; digit2<=TWO; digit3<=MIN; end
      16'd286: begin digit0<=SIX; digit1<=EIGHT; digit2<=TWO; digit3<=MIN; end
      16'd287: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=TWO; digit3<=MIN; end
      16'd288: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=TWO; digit3<=MIN; end
      16'd289: begin digit0<=NINE; digit1<=EIGHT; digit2<=TWO; digit3<=MIN; end
      16'd290: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=MIN; end
      16'd291: begin digit0<=ONE; digit1<=NINE; digit2<=TWO; digit3<=MIN; end
      16'd292: begin digit0<=ZERO; digit1<=NINE; digit2<=TWO; digit3<=MIN; end
      16'd293: begin digit0<=THREE; digit1<=NINE; digit2<=TWO; digit3<=MIN; end
      16'd294: begin digit0<=FOUR; digit1<=NINE; digit2<=TWO; digit3<=MIN; end
      16'd295: begin digit0<=FIVE; digit1<=NINE; digit2<=TWO; digit3<=MIN; end
      16'd296: begin digit0<=SIX; digit1<=NINE; digit2<=TWO; digit3<=MIN; end
      16'd297: begin digit0<=SEVEN; digit1<=NINE; digit2<=TWO; digit3<=MIN; end
      16'd298: begin digit0<=EIGHT; digit1<=NINE; digit2<=TWO; digit3<=MIN; end
      16'd299: begin digit0<=NINE; digit1<=NINE; digit2<=TWO; digit3<=MIN; end
	  16'd300: begin digit0<=ZERO; digit1<=ZERO; digit2<=THREE; digit3<=MIN; end
      16'd301: begin digit0<=ONE; digit1<=ZERO; digit2<=THREE; digit3<=MIN; end
      16'd302: begin digit0<=TWO; digit1<=ZERO; digit2<=THREE; digit3<=MIN; end
      16'd303: begin digit0<=THREE; digit1<=ZERO; digit2<=THREE; digit3<=MIN; end
      16'd304: begin digit0<=FOUR; digit1<=ZERO; digit2<=THREE; digit3<=MIN; end
      16'd305: begin digit0<=FIVE; digit1<=ZERO; digit2<=THREE; digit3<=MIN; end
      16'd306: begin digit0<=SIX; digit1<=ZERO; digit2<=THREE; digit3<=MIN; end
      16'd307: begin digit0<=SEVEN; digit1<=ZERO; digit2<=THREE; digit3<=MIN; end
      16'd308: begin digit0<=EIGHT; digit1<=ZERO; digit2<=THREE; digit3<=MIN; end
      16'd309: begin digit0<=NINE; digit1<=ZERO; digit2<=THREE; digit3<=MIN; end
      16'd310: begin digit0<=ZERO; digit1<=ONE; digit2<=THREE; digit3<=MIN; end
      16'd311: begin digit0<=ONE; digit1<=ONE; digit2<=THREE; digit3<=MIN; end
      16'd312: begin digit0<=TWO; digit1<=ONE; digit2<=THREE; digit3<=MIN; end
      16'd313: begin digit0<=THREE; digit1<=ONE; digit2<=THREE; digit3<=MIN; end
      16'd314: begin digit0<=FOUR; digit1<=ONE; digit2<=THREE; digit3<=MIN; end
      16'd315: begin digit0<=FIVE; digit1<=ONE; digit2<=THREE; digit3<=MIN; end
      16'd316: begin digit0<=SIX; digit1<=ONE; digit2<=THREE; digit3<=MIN; end
      16'd317: begin digit0<=SEVEN; digit1<=ONE; digit2<=THREE; digit3<=MIN; end
      16'd318: begin digit0<=EIGHT; digit1<=ONE; digit2<=THREE; digit3<=MIN; end
      16'd319: begin digit0<=NINE; digit1<=ONE; digit2<=THREE; digit3<=MIN; end
      16'd320: begin digit0<=ZERO; digit1<=TWO; digit2<=THREE; digit3<=MIN; end
      16'd321: begin digit0<=ONE; digit1<=TWO; digit2<=THREE; digit3<=MIN; end
      16'd322: begin digit0<=TWO; digit1<=TWO; digit2<=THREE; digit3<=MIN; end
      16'd323: begin digit0<=THREE; digit1<=TWO; digit2<=THREE; digit3<=MIN; end
      16'd324: begin digit0<=FOUR; digit1<=TWO; digit2<=THREE; digit3<=MIN; end
      16'd325: begin digit0<=FIVE; digit1<=TWO; digit2<=THREE; digit3<=MIN; end
      16'd326: begin digit0<=SIX; digit1<=TWO; digit2<=THREE; digit3<=MIN; end
      16'd327: begin digit0<=SEVEN; digit1<=TWO; digit2<=THREE; digit3<=MIN; end
      16'd328: begin digit0<=EIGHT; digit1<=TWO; digit2<=THREE; digit3<=MIN; end
      16'd329: begin digit0<=NINE; digit1<=TWO; digit2<=THREE; digit3<=MIN; end
      16'd330: begin digit0<=ZERO; digit1<=THREE; digit2<=THREE; digit3<=MIN; end
      16'd331: begin digit0<=ONE; digit1<=THREE; digit2<=THREE; digit3<=MIN; end
      16'd332: begin digit0<=TWO; digit1<=THREE; digit2<=THREE; digit3<=MIN; end
      16'd333: begin digit0<=THREE; digit1<=THREE; digit2<=THREE; digit3<=MIN; end
      16'd334: begin digit0<=FOUR; digit1<=THREE; digit2<=THREE; digit3<=MIN; end
      16'd335: begin digit0<=FIVE; digit1<=THREE; digit2<=THREE; digit3<=MIN; end
      16'd336: begin digit0<=SIX; digit1<=THREE; digit2<=THREE; digit3<=MIN; end
      16'd337: begin digit0<=SEVEN; digit1<=THREE; digit2<=THREE; digit3<=MIN; end
      16'd338: begin digit0<=EIGHT; digit1<=THREE; digit2<=THREE; digit3<=MIN; end
      16'd339: begin digit0<=NINE; digit1<=THREE; digit2<=THREE; digit3<=MIN; end
      16'd340: begin digit0<=ZERO; digit1<=FOUR; digit2<=THREE; digit3<=MIN; end
      16'd341: begin digit0<=ONE; digit1<=FOUR; digit2<=THREE; digit3<=MIN; end
      16'd342: begin digit0<=TWO; digit1<=FOUR; digit2<=THREE; digit3<=MIN; end
      16'd343: begin digit0<=THREE; digit1<=FOUR; digit2<=THREE; digit3<=MIN; end
      16'd344: begin digit0<=FOUR; digit1<=FOUR; digit2<=THREE; digit3<=MIN; end
      16'd345: begin digit0<=FIVE; digit1<=FOUR; digit2<=THREE; digit3<=MIN; end
      16'd346: begin digit0<=SIX; digit1<=FOUR; digit2<=THREE; digit3<=MIN; end
      16'd347: begin digit0<=SEVEN; digit1<=FOUR; digit2<=THREE; digit3<=MIN; end
      16'd348: begin digit0<=EIGHT; digit1<=FOUR; digit2<=THREE; digit3<=MIN; end
      16'd349: begin digit0<=NINE; digit1<=FOUR; digit2<=THREE; digit3<=MIN; end
      16'd350: begin digit0<=ZERO; digit1<=FIVE; digit2<=THREE; digit3<=MIN; end
      16'd351: begin digit0<=ONE; digit1<=FIVE; digit2<=THREE; digit3<=MIN; end
      16'd352: begin digit0<=TWO; digit1<=FIVE; digit2<=THREE; digit3<=MIN; end
      16'd353: begin digit0<=THREE; digit1<=FIVE; digit2<=THREE; digit3<=MIN; end
      16'd354: begin digit0<=FOUR; digit1<=FIVE; digit2<=THREE; digit3<=MIN; end
      16'd355: begin digit0<=FIVE; digit1<=FIVE; digit2<=THREE; digit3<=MIN; end
      16'd356: begin digit0<=SIX; digit1<=FIVE; digit2<=THREE; digit3<=MIN; end
      16'd357: begin digit0<=SEVEN; digit1<=FIVE; digit2<=THREE; digit3<=MIN; end
      16'd358: begin digit0<=EIGHT; digit1<=FIVE; digit2<=THREE; digit3<=MIN; end
      16'd359: begin digit0<=NINE; digit1<=FIVE; digit2<=THREE; digit3<=MIN; end
      16'd360: begin digit0<=ZERO; digit1<=SIX; digit2<=THREE; digit3<=MIN; end
      16'd361: begin digit0<=ONE; digit1<=SIX; digit2<=THREE; digit3<=MIN; end
      16'd362: begin digit0<=TWO; digit1<=SIX; digit2<=THREE; digit3<=MIN; end
      16'd363: begin digit0<=THREE; digit1<=SIX; digit2<=THREE; digit3<=MIN; end
      16'd364: begin digit0<=FOUR; digit1<=SIX; digit2<=THREE; digit3<=MIN; end
      16'd365: begin digit0<=FIVE; digit1<=SIX; digit2<=THREE; digit3<=MIN; end
      16'd366: begin digit0<=SIX; digit1<=SIX; digit2<=THREE; digit3<=MIN; end
      16'd367: begin digit0<=SEVEN; digit1<=SIX; digit2<=THREE; digit3<=MIN; end
      16'd368: begin digit0<=EIGHT; digit1<=SIX; digit2<=THREE; digit3<=MIN; end
      16'd369: begin digit0<=NINE; digit1<=SIX; digit2<=THREE; digit3<=MIN; end
      16'd370: begin digit0<=ZERO; digit1<=SEVEN; digit2<=THREE; digit3<=MIN; end
      16'd371: begin digit0<=ONE; digit1<=SEVEN; digit2<=THREE; digit3<=MIN; end
      16'd372: begin digit0<=TWO; digit1<=SEVEN; digit2<=THREE; digit3<=MIN; end
      16'd373: begin digit0<=THREE; digit1<=SEVEN; digit2<=THREE; digit3<=MIN; end
      16'd374: begin digit0<=FOUR; digit1<=SEVEN; digit2<=THREE; digit3<=MIN; end
      16'd375: begin digit0<=FIVE; digit1<=SEVEN; digit2<=THREE; digit3<=MIN; end
      16'd376: begin digit0<=SIX; digit1<=SEVEN; digit2<=THREE; digit3<=MIN; end
      16'd377: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=THREE; digit3<=MIN; end
      16'd378: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=THREE; digit3<=MIN; end
      16'd379: begin digit0<=NINE; digit1<=SEVEN; digit2<=THREE; digit3<=MIN; end
      16'd380: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=MIN; end
      16'd381: begin digit0<=ONE; digit1<=EIGHT; digit2<=THREE; digit3<=MIN; end
      16'd382: begin digit0<=ZERO; digit1<=EIGHT; digit2<=THREE; digit3<=MIN; end
      16'd383: begin digit0<=THREE; digit1<=EIGHT; digit2<=THREE; digit3<=MIN; end
      16'd384: begin digit0<=FOUR; digit1<=EIGHT; digit2<=THREE; digit3<=MIN; end
      16'd385: begin digit0<=FIVE; digit1<=EIGHT; digit2<=THREE; digit3<=MIN; end
      16'd386: begin digit0<=SIX; digit1<=EIGHT; digit2<=THREE; digit3<=MIN; end
      16'd387: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=THREE; digit3<=MIN; end
      16'd388: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=THREE; digit3<=MIN; end
      16'd389: begin digit0<=NINE; digit1<=EIGHT; digit2<=THREE; digit3<=MIN; end
      16'd390: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=MIN; end
      16'd391: begin digit0<=ONE; digit1<=NINE; digit2<=THREE; digit3<=MIN; end
      16'd392: begin digit0<=ZERO; digit1<=NINE; digit2<=THREE; digit3<=MIN; end
      16'd393: begin digit0<=THREE; digit1<=NINE; digit2<=THREE; digit3<=MIN; end
      16'd394: begin digit0<=FOUR; digit1<=NINE; digit2<=THREE; digit3<=MIN; end
      16'd395: begin digit0<=FIVE; digit1<=NINE; digit2<=THREE; digit3<=MIN; end
      16'd396: begin digit0<=SIX; digit1<=NINE; digit2<=THREE; digit3<=MIN; end
      16'd397: begin digit0<=SEVEN; digit1<=NINE; digit2<=THREE; digit3<=MIN; end
      16'd398: begin digit0<=EIGHT; digit1<=NINE; digit2<=THREE; digit3<=MIN; end
      16'd399: begin digit0<=NINE; digit1<=NINE; digit2<=THREE; digit3<=MIN; end
	  16'd400: begin digit0<=ZERO; digit1<=ZERO; digit2<=FOUR; digit3<=MIN; end
      16'd401: begin digit0<=ONE; digit1<=ZERO; digit2<=FOUR; digit3<=MIN; end
      16'd402: begin digit0<=TWO; digit1<=ZERO; digit2<=FOUR; digit3<=MIN; end
      16'd403: begin digit0<=THREE; digit1<=ZERO; digit2<=FOUR; digit3<=MIN; end
      16'd404: begin digit0<=FOUR; digit1<=ZERO; digit2<=FOUR; digit3<=MIN; end
      16'd405: begin digit0<=FIVE; digit1<=ZERO; digit2<=FOUR; digit3<=MIN; end
      16'd406: begin digit0<=SIX; digit1<=ZERO; digit2<=FOUR; digit3<=MIN; end
      16'd407: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FOUR; digit3<=MIN; end
      16'd408: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FOUR; digit3<=MIN; end
      16'd409: begin digit0<=NINE; digit1<=ZERO; digit2<=FOUR; digit3<=MIN; end
      16'd410: begin digit0<=ZERO; digit1<=ONE; digit2<=FOUR; digit3<=MIN; end
      16'd411: begin digit0<=ONE; digit1<=ONE; digit2<=FOUR; digit3<=MIN; end
      16'd412: begin digit0<=TWO; digit1<=ONE; digit2<=FOUR; digit3<=MIN; end
      16'd413: begin digit0<=THREE; digit1<=ONE; digit2<=FOUR; digit3<=MIN; end
      16'd414: begin digit0<=FOUR; digit1<=ONE; digit2<=FOUR; digit3<=MIN; end
      16'd415: begin digit0<=FIVE; digit1<=ONE; digit2<=FOUR; digit3<=MIN; end
      16'd416: begin digit0<=SIX; digit1<=ONE; digit2<=FOUR; digit3<=MIN; end
      16'd417: begin digit0<=SEVEN; digit1<=ONE; digit2<=FOUR; digit3<=MIN; end
      16'd418: begin digit0<=EIGHT; digit1<=ONE; digit2<=FOUR; digit3<=MIN; end
      16'd419: begin digit0<=NINE; digit1<=ONE; digit2<=FOUR; digit3<=MIN; end
      16'd420: begin digit0<=ZERO; digit1<=TWO; digit2<=FOUR; digit3<=MIN; end
      16'd421: begin digit0<=ONE; digit1<=TWO; digit2<=FOUR; digit3<=MIN; end
      16'd422: begin digit0<=TWO; digit1<=TWO; digit2<=FOUR; digit3<=MIN; end
      16'd423: begin digit0<=THREE; digit1<=TWO; digit2<=FOUR; digit3<=MIN; end
      16'd424: begin digit0<=FOUR; digit1<=TWO; digit2<=FOUR; digit3<=MIN; end
      16'd425: begin digit0<=FIVE; digit1<=TWO; digit2<=FOUR; digit3<=MIN; end
      16'd426: begin digit0<=SIX; digit1<=TWO; digit2<=FOUR; digit3<=MIN; end
      16'd427: begin digit0<=SEVEN; digit1<=TWO; digit2<=FOUR; digit3<=MIN; end
      16'd428: begin digit0<=EIGHT; digit1<=TWO; digit2<=FOUR; digit3<=MIN; end
      16'd429: begin digit0<=NINE; digit1<=TWO; digit2<=FOUR; digit3<=MIN; end
      16'd430: begin digit0<=ZERO; digit1<=THREE; digit2<=FOUR; digit3<=MIN; end
      16'd431: begin digit0<=ONE; digit1<=THREE; digit2<=FOUR; digit3<=MIN; end
      16'd432: begin digit0<=TWO; digit1<=THREE; digit2<=FOUR; digit3<=MIN; end
      16'd433: begin digit0<=THREE; digit1<=THREE; digit2<=FOUR; digit3<=MIN; end
      16'd434: begin digit0<=FOUR; digit1<=THREE; digit2<=FOUR; digit3<=MIN; end
      16'd435: begin digit0<=FIVE; digit1<=THREE; digit2<=FOUR; digit3<=MIN; end
      16'd436: begin digit0<=SIX; digit1<=THREE; digit2<=FOUR; digit3<=MIN; end
      16'd437: begin digit0<=SEVEN; digit1<=THREE; digit2<=FOUR; digit3<=MIN; end
      16'd438: begin digit0<=EIGHT; digit1<=THREE; digit2<=FOUR; digit3<=MIN; end
      16'd439: begin digit0<=NINE; digit1<=THREE; digit2<=FOUR; digit3<=MIN; end
      16'd440: begin digit0<=ZERO; digit1<=FOUR; digit2<=FOUR; digit3<=MIN; end
      16'd441: begin digit0<=ONE; digit1<=FOUR; digit2<=FOUR; digit3<=MIN; end
      16'd442: begin digit0<=TWO; digit1<=FOUR; digit2<=FOUR; digit3<=MIN; end
      16'd443: begin digit0<=THREE; digit1<=FOUR; digit2<=FOUR; digit3<=MIN; end
      16'd444: begin digit0<=FOUR; digit1<=FOUR; digit2<=FOUR; digit3<=MIN; end
      16'd445: begin digit0<=FIVE; digit1<=FOUR; digit2<=FOUR; digit3<=MIN; end
      16'd446: begin digit0<=SIX; digit1<=FOUR; digit2<=FOUR; digit3<=MIN; end
      16'd447: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FOUR; digit3<=MIN; end
      16'd448: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FOUR; digit3<=MIN; end
      16'd449: begin digit0<=NINE; digit1<=FOUR; digit2<=FOUR; digit3<=MIN; end
      16'd450: begin digit0<=ZERO; digit1<=FIVE; digit2<=FOUR; digit3<=MIN; end
      16'd451: begin digit0<=ONE; digit1<=FIVE; digit2<=FOUR; digit3<=MIN; end
      16'd452: begin digit0<=TWO; digit1<=FIVE; digit2<=FOUR; digit3<=MIN; end
      16'd453: begin digit0<=THREE; digit1<=FIVE; digit2<=FOUR; digit3<=MIN; end
      16'd454: begin digit0<=FOUR; digit1<=FIVE; digit2<=FOUR; digit3<=MIN; end
      16'd455: begin digit0<=FIVE; digit1<=FIVE; digit2<=FOUR; digit3<=MIN; end
      16'd456: begin digit0<=SIX; digit1<=FIVE; digit2<=FOUR; digit3<=MIN; end
      16'd457: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FOUR; digit3<=MIN; end
      16'd458: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FOUR; digit3<=MIN; end
      16'd459: begin digit0<=NINE; digit1<=FIVE; digit2<=FOUR; digit3<=MIN; end
      16'd460: begin digit0<=ZERO; digit1<=SIX; digit2<=FOUR; digit3<=MIN; end
      16'd461: begin digit0<=ONE; digit1<=SIX; digit2<=FOUR; digit3<=MIN; end
      16'd462: begin digit0<=TWO; digit1<=SIX; digit2<=FOUR; digit3<=MIN; end
      16'd463: begin digit0<=THREE; digit1<=SIX; digit2<=FOUR; digit3<=MIN; end
      16'd464: begin digit0<=FOUR; digit1<=SIX; digit2<=FOUR; digit3<=MIN; end
      16'd465: begin digit0<=FIVE; digit1<=SIX; digit2<=FOUR; digit3<=MIN; end
      16'd466: begin digit0<=SIX; digit1<=SIX; digit2<=FOUR; digit3<=MIN; end
      16'd467: begin digit0<=SEVEN; digit1<=SIX; digit2<=FOUR; digit3<=MIN; end
      16'd468: begin digit0<=EIGHT; digit1<=SIX; digit2<=FOUR; digit3<=MIN; end
      16'd469: begin digit0<=NINE; digit1<=SIX; digit2<=FOUR; digit3<=MIN; end
      16'd470: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FOUR; digit3<=MIN; end
      16'd471: begin digit0<=ONE; digit1<=SEVEN; digit2<=FOUR; digit3<=MIN; end
      16'd472: begin digit0<=TWO; digit1<=SEVEN; digit2<=FOUR; digit3<=MIN; end
      16'd473: begin digit0<=THREE; digit1<=SEVEN; digit2<=FOUR; digit3<=MIN; end
      16'd474: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FOUR; digit3<=MIN; end
      16'd475: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FOUR; digit3<=MIN; end
      16'd476: begin digit0<=SIX; digit1<=SEVEN; digit2<=FOUR; digit3<=MIN; end
      16'd477: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FOUR; digit3<=MIN; end
      16'd478: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FOUR; digit3<=MIN; end
      16'd479: begin digit0<=NINE; digit1<=SEVEN; digit2<=FOUR; digit3<=MIN; end
      16'd480: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=MIN; end
      16'd481: begin digit0<=ONE; digit1<=EIGHT; digit2<=FOUR; digit3<=MIN; end
      16'd482: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FOUR; digit3<=MIN; end
      16'd483: begin digit0<=THREE; digit1<=EIGHT; digit2<=FOUR; digit3<=MIN; end
      16'd484: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FOUR; digit3<=MIN; end
      16'd485: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FOUR; digit3<=MIN; end
      16'd486: begin digit0<=SIX; digit1<=EIGHT; digit2<=FOUR; digit3<=MIN; end
      16'd487: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FOUR; digit3<=MIN; end
      16'd488: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FOUR; digit3<=MIN; end
      16'd489: begin digit0<=NINE; digit1<=EIGHT; digit2<=FOUR; digit3<=MIN; end
      16'd490: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=MIN; end
      16'd491: begin digit0<=ONE; digit1<=NINE; digit2<=FOUR; digit3<=MIN; end
      16'd492: begin digit0<=ZERO; digit1<=NINE; digit2<=FOUR; digit3<=MIN; end
      16'd493: begin digit0<=THREE; digit1<=NINE; digit2<=FOUR; digit3<=MIN; end
      16'd494: begin digit0<=FOUR; digit1<=NINE; digit2<=FOUR; digit3<=MIN; end
      16'd495: begin digit0<=FIVE; digit1<=NINE; digit2<=FOUR; digit3<=MIN; end
      16'd496: begin digit0<=SIX; digit1<=NINE; digit2<=FOUR; digit3<=MIN; end
      16'd497: begin digit0<=SEVEN; digit1<=NINE; digit2<=FOUR; digit3<=MIN; end
      16'd498: begin digit0<=EIGHT; digit1<=NINE; digit2<=FOUR; digit3<=MIN; end
      16'd499: begin digit0<=NINE; digit1<=NINE; digit2<=FOUR; digit3<=MIN; end
	  16'd500: begin digit0<=ZERO; digit1<=ZERO; digit2<=FIVE; digit3<=MIN; end
      16'd501: begin digit0<=ONE; digit1<=ZERO; digit2<=FIVE; digit3<=MIN; end
      16'd502: begin digit0<=TWO; digit1<=ZERO; digit2<=FIVE; digit3<=MIN; end
      16'd503: begin digit0<=THREE; digit1<=ZERO; digit2<=FIVE; digit3<=MIN; end
      16'd504: begin digit0<=FOUR; digit1<=ZERO; digit2<=FIVE; digit3<=MIN; end
      16'd505: begin digit0<=FIVE; digit1<=ZERO; digit2<=FIVE; digit3<=MIN; end
      16'd506: begin digit0<=SIX; digit1<=ZERO; digit2<=FIVE; digit3<=MIN; end
      16'd507: begin digit0<=SEVEN; digit1<=ZERO; digit2<=FIVE; digit3<=MIN; end
      16'd508: begin digit0<=EIGHT; digit1<=ZERO; digit2<=FIVE; digit3<=MIN; end
      16'd509: begin digit0<=NINE; digit1<=ZERO; digit2<=FIVE; digit3<=MIN; end
      16'd510: begin digit0<=ZERO; digit1<=ONE; digit2<=FIVE; digit3<=MIN; end
      16'd511: begin digit0<=ONE; digit1<=ONE; digit2<=FIVE; digit3<=MIN; end
      16'd512: begin digit0<=TWO; digit1<=ONE; digit2<=FIVE; digit3<=MIN; end
      16'd513: begin digit0<=THREE; digit1<=ONE; digit2<=FIVE; digit3<=MIN; end
      16'd514: begin digit0<=FOUR; digit1<=ONE; digit2<=FIVE; digit3<=MIN; end
      16'd515: begin digit0<=FIVE; digit1<=ONE; digit2<=FIVE; digit3<=MIN; end
      16'd516: begin digit0<=SIX; digit1<=ONE; digit2<=FIVE; digit3<=MIN; end
      16'd517: begin digit0<=SEVEN; digit1<=ONE; digit2<=FIVE; digit3<=MIN; end
      16'd518: begin digit0<=EIGHT; digit1<=ONE; digit2<=FIVE; digit3<=MIN; end
      16'd519: begin digit0<=NINE; digit1<=ONE; digit2<=FIVE; digit3<=MIN; end
      16'd520: begin digit0<=ZERO; digit1<=TWO; digit2<=FIVE; digit3<=MIN; end
      16'd521: begin digit0<=ONE; digit1<=TWO; digit2<=FIVE; digit3<=MIN; end
      16'd522: begin digit0<=TWO; digit1<=TWO; digit2<=FIVE; digit3<=MIN; end
      16'd523: begin digit0<=THREE; digit1<=TWO; digit2<=FIVE; digit3<=MIN; end
      16'd524: begin digit0<=FOUR; digit1<=TWO; digit2<=FIVE; digit3<=MIN; end
      16'd525: begin digit0<=FIVE; digit1<=TWO; digit2<=FIVE; digit3<=MIN; end
      16'd526: begin digit0<=SIX; digit1<=TWO; digit2<=FIVE; digit3<=MIN; end
      16'd527: begin digit0<=SEVEN; digit1<=TWO; digit2<=FIVE; digit3<=MIN; end
      16'd528: begin digit0<=EIGHT; digit1<=TWO; digit2<=FIVE; digit3<=MIN; end
      16'd529: begin digit0<=NINE; digit1<=TWO; digit2<=FIVE; digit3<=MIN; end
      16'd530: begin digit0<=ZERO; digit1<=THREE; digit2<=FIVE; digit3<=MIN; end
      16'd531: begin digit0<=ONE; digit1<=THREE; digit2<=FIVE; digit3<=MIN; end
      16'd532: begin digit0<=TWO; digit1<=THREE; digit2<=FIVE; digit3<=MIN; end
      16'd533: begin digit0<=THREE; digit1<=THREE; digit2<=FIVE; digit3<=MIN; end
      16'd534: begin digit0<=FOUR; digit1<=THREE; digit2<=FIVE; digit3<=MIN; end
      16'd535: begin digit0<=FIVE; digit1<=THREE; digit2<=FIVE; digit3<=MIN; end
      16'd536: begin digit0<=SIX; digit1<=THREE; digit2<=FIVE; digit3<=MIN; end
      16'd537: begin digit0<=SEVEN; digit1<=THREE; digit2<=FIVE; digit3<=MIN; end
      16'd538: begin digit0<=EIGHT; digit1<=THREE; digit2<=FIVE; digit3<=MIN; end
      16'd539: begin digit0<=NINE; digit1<=THREE; digit2<=FIVE; digit3<=MIN; end
      16'd540: begin digit0<=ZERO; digit1<=FOUR; digit2<=FIVE; digit3<=MIN; end
      16'd541: begin digit0<=ONE; digit1<=FOUR; digit2<=FIVE; digit3<=MIN; end
      16'd542: begin digit0<=TWO; digit1<=FOUR; digit2<=FIVE; digit3<=MIN; end
      16'd543: begin digit0<=THREE; digit1<=FOUR; digit2<=FIVE; digit3<=MIN; end
      16'd544: begin digit0<=FOUR; digit1<=FOUR; digit2<=FIVE; digit3<=MIN; end
      16'd545: begin digit0<=FIVE; digit1<=FOUR; digit2<=FIVE; digit3<=MIN; end
      16'd546: begin digit0<=SIX; digit1<=FOUR; digit2<=FIVE; digit3<=MIN; end
      16'd547: begin digit0<=SEVEN; digit1<=FOUR; digit2<=FIVE; digit3<=MIN; end
      16'd548: begin digit0<=EIGHT; digit1<=FOUR; digit2<=FIVE; digit3<=MIN; end
      16'd549: begin digit0<=NINE; digit1<=FOUR; digit2<=FIVE; digit3<=MIN; end
      16'd550: begin digit0<=ZERO; digit1<=FIVE; digit2<=FIVE; digit3<=MIN; end
      16'd551: begin digit0<=ONE; digit1<=FIVE; digit2<=FIVE; digit3<=MIN; end
      16'd552: begin digit0<=TWO; digit1<=FIVE; digit2<=FIVE; digit3<=MIN; end
      16'd553: begin digit0<=THREE; digit1<=FIVE; digit2<=FIVE; digit3<=MIN; end
      16'd554: begin digit0<=FOUR; digit1<=FIVE; digit2<=FIVE; digit3<=MIN; end
      16'd555: begin digit0<=FIVE; digit1<=FIVE; digit2<=FIVE; digit3<=MIN; end
      16'd556: begin digit0<=SIX; digit1<=FIVE; digit2<=FIVE; digit3<=MIN; end
      16'd557: begin digit0<=SEVEN; digit1<=FIVE; digit2<=FIVE; digit3<=MIN; end
      16'd558: begin digit0<=EIGHT; digit1<=FIVE; digit2<=FIVE; digit3<=MIN; end
      16'd559: begin digit0<=NINE; digit1<=FIVE; digit2<=FIVE; digit3<=MIN; end
      16'd560: begin digit0<=ZERO; digit1<=SIX; digit2<=FIVE; digit3<=MIN; end
      16'd561: begin digit0<=ONE; digit1<=SIX; digit2<=FIVE; digit3<=MIN; end
      16'd562: begin digit0<=TWO; digit1<=SIX; digit2<=FIVE; digit3<=MIN; end
      16'd563: begin digit0<=THREE; digit1<=SIX; digit2<=FIVE; digit3<=MIN; end
      16'd564: begin digit0<=FOUR; digit1<=SIX; digit2<=FIVE; digit3<=MIN; end
      16'd565: begin digit0<=FIVE; digit1<=SIX; digit2<=FIVE; digit3<=MIN; end
      16'd566: begin digit0<=SIX; digit1<=SIX; digit2<=FIVE; digit3<=MIN; end
      16'd567: begin digit0<=SEVEN; digit1<=SIX; digit2<=FIVE; digit3<=MIN; end
      16'd568: begin digit0<=EIGHT; digit1<=SIX; digit2<=FIVE; digit3<=MIN; end
      16'd569: begin digit0<=NINE; digit1<=SIX; digit2<=FIVE; digit3<=MIN; end
      16'd570: begin digit0<=ZERO; digit1<=SEVEN; digit2<=FIVE; digit3<=MIN; end
      16'd571: begin digit0<=ONE; digit1<=SEVEN; digit2<=FIVE; digit3<=MIN; end
      16'd572: begin digit0<=TWO; digit1<=SEVEN; digit2<=FIVE; digit3<=MIN; end
      16'd573: begin digit0<=THREE; digit1<=SEVEN; digit2<=FIVE; digit3<=MIN; end
      16'd574: begin digit0<=FOUR; digit1<=SEVEN; digit2<=FIVE; digit3<=MIN; end
      16'd575: begin digit0<=FIVE; digit1<=SEVEN; digit2<=FIVE; digit3<=MIN; end
      16'd576: begin digit0<=SIX; digit1<=SEVEN; digit2<=FIVE; digit3<=MIN; end
      16'd577: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=FIVE; digit3<=MIN; end
      16'd578: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=FIVE; digit3<=MIN; end
      16'd579: begin digit0<=NINE; digit1<=SEVEN; digit2<=FIVE; digit3<=MIN; end
      16'd580: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=MIN; end
      16'd581: begin digit0<=ONE; digit1<=EIGHT; digit2<=FIVE; digit3<=MIN; end
      16'd582: begin digit0<=ZERO; digit1<=EIGHT; digit2<=FIVE; digit3<=MIN; end
      16'd583: begin digit0<=THREE; digit1<=EIGHT; digit2<=FIVE; digit3<=MIN; end
      16'd584: begin digit0<=FOUR; digit1<=EIGHT; digit2<=FIVE; digit3<=MIN; end
      16'd585: begin digit0<=FIVE; digit1<=EIGHT; digit2<=FIVE; digit3<=MIN; end
      16'd586: begin digit0<=SIX; digit1<=EIGHT; digit2<=FIVE; digit3<=MIN; end
      16'd587: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=FIVE; digit3<=MIN; end
      16'd588: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=FIVE; digit3<=MIN; end
      16'd589: begin digit0<=NINE; digit1<=EIGHT; digit2<=FIVE; digit3<=MIN; end
      16'd590: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=MIN; end
      16'd591: begin digit0<=ONE; digit1<=NINE; digit2<=FIVE; digit3<=MIN; end
      16'd592: begin digit0<=ZERO; digit1<=NINE; digit2<=FIVE; digit3<=MIN; end
      16'd593: begin digit0<=THREE; digit1<=NINE; digit2<=FIVE; digit3<=MIN; end
      16'd594: begin digit0<=FOUR; digit1<=NINE; digit2<=FIVE; digit3<=MIN; end
      16'd595: begin digit0<=FIVE; digit1<=NINE; digit2<=FIVE; digit3<=MIN; end
      16'd596: begin digit0<=SIX; digit1<=NINE; digit2<=FIVE; digit3<=MIN; end
      16'd597: begin digit0<=SEVEN; digit1<=NINE; digit2<=FIVE; digit3<=MIN; end
      16'd598: begin digit0<=EIGHT; digit1<=NINE; digit2<=FIVE; digit3<=MIN; end
      16'd599: begin digit0<=NINE; digit1<=NINE; digit2<=FIVE; digit3<=MIN; end
	  16'd600: begin digit0<=ZERO; digit1<=ZERO; digit2<=SIX; digit3<=MIN; end
      16'd601: begin digit0<=ONE; digit1<=ZERO; digit2<=SIX; digit3<=MIN; end
      16'd602: begin digit0<=TWO; digit1<=ZERO; digit2<=SIX; digit3<=MIN; end
      16'd603: begin digit0<=THREE; digit1<=ZERO; digit2<=SIX; digit3<=MIN; end
      16'd604: begin digit0<=FOUR; digit1<=ZERO; digit2<=SIX; digit3<=MIN; end
      16'd605: begin digit0<=FIVE; digit1<=ZERO; digit2<=SIX; digit3<=MIN; end
      16'd606: begin digit0<=SIX; digit1<=ZERO; digit2<=SIX; digit3<=MIN; end
      16'd607: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SIX; digit3<=MIN; end
      16'd608: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SIX; digit3<=MIN; end
      16'd609: begin digit0<=NINE; digit1<=ZERO; digit2<=SIX; digit3<=MIN; end
      16'd610: begin digit0<=ZERO; digit1<=ONE; digit2<=SIX; digit3<=MIN; end
      16'd611: begin digit0<=ONE; digit1<=ONE; digit2<=SIX; digit3<=MIN; end
      16'd612: begin digit0<=TWO; digit1<=ONE; digit2<=SIX; digit3<=MIN; end
      16'd613: begin digit0<=THREE; digit1<=ONE; digit2<=SIX; digit3<=MIN; end
      16'd614: begin digit0<=FOUR; digit1<=ONE; digit2<=SIX; digit3<=MIN; end
      16'd615: begin digit0<=FIVE; digit1<=ONE; digit2<=SIX; digit3<=MIN; end
      16'd616: begin digit0<=SIX; digit1<=ONE; digit2<=SIX; digit3<=MIN; end
      16'd617: begin digit0<=SEVEN; digit1<=ONE; digit2<=SIX; digit3<=MIN; end
      16'd618: begin digit0<=EIGHT; digit1<=ONE; digit2<=SIX; digit3<=MIN; end
      16'd619: begin digit0<=NINE; digit1<=ONE; digit2<=SIX; digit3<=MIN; end
      16'd620: begin digit0<=ZERO; digit1<=TWO; digit2<=SIX; digit3<=MIN; end
      16'd621: begin digit0<=ONE; digit1<=TWO; digit2<=SIX; digit3<=MIN; end
      16'd622: begin digit0<=TWO; digit1<=TWO; digit2<=SIX; digit3<=MIN; end
      16'd623: begin digit0<=THREE; digit1<=TWO; digit2<=SIX; digit3<=MIN; end
      16'd624: begin digit0<=FOUR; digit1<=TWO; digit2<=SIX; digit3<=MIN; end
      16'd625: begin digit0<=FIVE; digit1<=TWO; digit2<=SIX; digit3<=MIN; end
      16'd626: begin digit0<=SIX; digit1<=TWO; digit2<=SIX; digit3<=MIN; end
      16'd627: begin digit0<=SEVEN; digit1<=TWO; digit2<=SIX; digit3<=MIN; end
      16'd628: begin digit0<=EIGHT; digit1<=TWO; digit2<=SIX; digit3<=MIN; end
      16'd629: begin digit0<=NINE; digit1<=TWO; digit2<=SIX; digit3<=MIN; end
      16'd630: begin digit0<=ZERO; digit1<=THREE; digit2<=SIX; digit3<=MIN; end
      16'd631: begin digit0<=ONE; digit1<=THREE; digit2<=SIX; digit3<=MIN; end
      16'd632: begin digit0<=TWO; digit1<=THREE; digit2<=SIX; digit3<=MIN; end
      16'd633: begin digit0<=THREE; digit1<=THREE; digit2<=SIX; digit3<=MIN; end
      16'd634: begin digit0<=FOUR; digit1<=THREE; digit2<=SIX; digit3<=MIN; end
      16'd635: begin digit0<=FIVE; digit1<=THREE; digit2<=SIX; digit3<=MIN; end
      16'd636: begin digit0<=SIX; digit1<=THREE; digit2<=SIX; digit3<=MIN; end
      16'd637: begin digit0<=SEVEN; digit1<=THREE; digit2<=SIX; digit3<=MIN; end
      16'd638: begin digit0<=EIGHT; digit1<=THREE; digit2<=SIX; digit3<=MIN; end
      16'd639: begin digit0<=NINE; digit1<=THREE; digit2<=SIX; digit3<=MIN; end
      16'd640: begin digit0<=ZERO; digit1<=FOUR; digit2<=SIX; digit3<=MIN; end
      16'd641: begin digit0<=ONE; digit1<=FOUR; digit2<=SIX; digit3<=MIN; end
      16'd642: begin digit0<=TWO; digit1<=FOUR; digit2<=SIX; digit3<=MIN; end
      16'd643: begin digit0<=THREE; digit1<=FOUR; digit2<=SIX; digit3<=MIN; end
      16'd644: begin digit0<=FOUR; digit1<=FOUR; digit2<=SIX; digit3<=MIN; end
      16'd645: begin digit0<=FIVE; digit1<=FOUR; digit2<=SIX; digit3<=MIN; end
      16'd646: begin digit0<=SIX; digit1<=FOUR; digit2<=SIX; digit3<=MIN; end
      16'd647: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SIX; digit3<=MIN; end
      16'd648: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SIX; digit3<=MIN; end
      16'd649: begin digit0<=NINE; digit1<=FOUR; digit2<=SIX; digit3<=MIN; end
      16'd650: begin digit0<=ZERO; digit1<=FIVE; digit2<=SIX; digit3<=MIN; end
      16'd651: begin digit0<=ONE; digit1<=FIVE; digit2<=SIX; digit3<=MIN; end
      16'd652: begin digit0<=TWO; digit1<=FIVE; digit2<=SIX; digit3<=MIN; end
      16'd653: begin digit0<=THREE; digit1<=FIVE; digit2<=SIX; digit3<=MIN; end
      16'd654: begin digit0<=FOUR; digit1<=FIVE; digit2<=SIX; digit3<=MIN; end
      16'd655: begin digit0<=FIVE; digit1<=FIVE; digit2<=SIX; digit3<=MIN; end
      16'd656: begin digit0<=SIX; digit1<=FIVE; digit2<=SIX; digit3<=MIN; end
      16'd657: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SIX; digit3<=MIN; end
      16'd658: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SIX; digit3<=MIN; end
      16'd659: begin digit0<=NINE; digit1<=FIVE; digit2<=SIX; digit3<=MIN; end
      16'd660: begin digit0<=ZERO; digit1<=SIX; digit2<=SIX; digit3<=MIN; end
      16'd661: begin digit0<=ONE; digit1<=SIX; digit2<=SIX; digit3<=MIN; end
      16'd662: begin digit0<=TWO; digit1<=SIX; digit2<=SIX; digit3<=MIN; end
      16'd663: begin digit0<=THREE; digit1<=SIX; digit2<=SIX; digit3<=MIN; end
      16'd664: begin digit0<=FOUR; digit1<=SIX; digit2<=SIX; digit3<=MIN; end
      16'd665: begin digit0<=FIVE; digit1<=SIX; digit2<=SIX; digit3<=MIN; end
      16'd666: begin digit0<=SIX; digit1<=SIX; digit2<=SIX; digit3<=MIN; end
      16'd667: begin digit0<=SEVEN; digit1<=SIX; digit2<=SIX; digit3<=MIN; end
      16'd668: begin digit0<=EIGHT; digit1<=SIX; digit2<=SIX; digit3<=MIN; end
      16'd669: begin digit0<=NINE; digit1<=SIX; digit2<=SIX; digit3<=MIN; end
      16'd670: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SIX; digit3<=MIN; end
      16'd671: begin digit0<=ONE; digit1<=SEVEN; digit2<=SIX; digit3<=MIN; end
      16'd672: begin digit0<=TWO; digit1<=SEVEN; digit2<=SIX; digit3<=MIN; end
      16'd673: begin digit0<=THREE; digit1<=SEVEN; digit2<=SIX; digit3<=MIN; end
      16'd674: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SIX; digit3<=MIN; end
      16'd675: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SIX; digit3<=MIN; end
      16'd676: begin digit0<=SIX; digit1<=SEVEN; digit2<=SIX; digit3<=MIN; end
      16'd677: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SIX; digit3<=MIN; end
      16'd678: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SIX; digit3<=MIN; end
      16'd679: begin digit0<=NINE; digit1<=SEVEN; digit2<=SIX; digit3<=MIN; end
      16'd680: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=MIN; end
      16'd681: begin digit0<=ONE; digit1<=EIGHT; digit2<=SIX; digit3<=MIN; end
      16'd682: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SIX; digit3<=MIN; end
      16'd683: begin digit0<=THREE; digit1<=EIGHT; digit2<=SIX; digit3<=MIN; end
      16'd684: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SIX; digit3<=MIN; end
      16'd685: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SIX; digit3<=MIN; end
      16'd686: begin digit0<=SIX; digit1<=EIGHT; digit2<=SIX; digit3<=MIN; end
      16'd687: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SIX; digit3<=MIN; end
      16'd688: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SIX; digit3<=MIN; end
      16'd689: begin digit0<=NINE; digit1<=EIGHT; digit2<=SIX; digit3<=MIN; end
      16'd690: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=MIN; end
      16'd691: begin digit0<=ONE; digit1<=NINE; digit2<=SIX; digit3<=MIN; end
      16'd692: begin digit0<=ZERO; digit1<=NINE; digit2<=SIX; digit3<=MIN; end
      16'd693: begin digit0<=THREE; digit1<=NINE; digit2<=SIX; digit3<=MIN; end
      16'd694: begin digit0<=FOUR; digit1<=NINE; digit2<=SIX; digit3<=MIN; end
      16'd695: begin digit0<=FIVE; digit1<=NINE; digit2<=SIX; digit3<=MIN; end
      16'd696: begin digit0<=SIX; digit1<=NINE; digit2<=SIX; digit3<=MIN; end
      16'd697: begin digit0<=SEVEN; digit1<=NINE; digit2<=SIX; digit3<=MIN; end
      16'd698: begin digit0<=EIGHT; digit1<=NINE; digit2<=SIX; digit3<=MIN; end
      16'd699: begin digit0<=NINE; digit1<=NINE; digit2<=SIX; digit3<=MIN; end
	  16'd700: begin digit0<=ZERO; digit1<=ZERO; digit2<=SEVEN; digit3<=MIN; end
      16'd701: begin digit0<=ONE; digit1<=ZERO; digit2<=SEVEN; digit3<=MIN; end
      16'd702: begin digit0<=TWO; digit1<=ZERO; digit2<=SEVEN; digit3<=MIN; end
      16'd703: begin digit0<=THREE; digit1<=ZERO; digit2<=SEVEN; digit3<=MIN; end
      16'd704: begin digit0<=FOUR; digit1<=ZERO; digit2<=SEVEN; digit3<=MIN; end
      16'd705: begin digit0<=FIVE; digit1<=ZERO; digit2<=SEVEN; digit3<=MIN; end
      16'd706: begin digit0<=SIX; digit1<=ZERO; digit2<=SEVEN; digit3<=MIN; end
      16'd707: begin digit0<=SEVEN; digit1<=ZERO; digit2<=SEVEN; digit3<=MIN; end
      16'd708: begin digit0<=EIGHT; digit1<=ZERO; digit2<=SEVEN; digit3<=MIN; end
      16'd709: begin digit0<=NINE; digit1<=ZERO; digit2<=SEVEN; digit3<=MIN; end
      16'd710: begin digit0<=ZERO; digit1<=ONE; digit2<=SEVEN; digit3<=MIN; end
      16'd711: begin digit0<=ONE; digit1<=ONE; digit2<=SEVEN; digit3<=MIN; end
      16'd712: begin digit0<=TWO; digit1<=ONE; digit2<=SEVEN; digit3<=MIN; end
      16'd713: begin digit0<=THREE; digit1<=ONE; digit2<=SEVEN; digit3<=MIN; end
      16'd714: begin digit0<=FOUR; digit1<=ONE; digit2<=SEVEN; digit3<=MIN; end
      16'd715: begin digit0<=FIVE; digit1<=ONE; digit2<=SEVEN; digit3<=MIN; end
      16'd716: begin digit0<=SIX; digit1<=ONE; digit2<=SEVEN; digit3<=MIN; end
      16'd717: begin digit0<=SEVEN; digit1<=ONE; digit2<=SEVEN; digit3<=MIN; end
      16'd718: begin digit0<=EIGHT; digit1<=ONE; digit2<=SEVEN; digit3<=MIN; end
      16'd719: begin digit0<=NINE; digit1<=ONE; digit2<=SEVEN; digit3<=MIN; end
      16'd720: begin digit0<=ZERO; digit1<=TWO; digit2<=SEVEN; digit3<=MIN; end
      16'd721: begin digit0<=ONE; digit1<=TWO; digit2<=SEVEN; digit3<=MIN; end
      16'd722: begin digit0<=TWO; digit1<=TWO; digit2<=SEVEN; digit3<=MIN; end
      16'd723: begin digit0<=THREE; digit1<=TWO; digit2<=SEVEN; digit3<=MIN; end
      16'd724: begin digit0<=FOUR; digit1<=TWO; digit2<=SEVEN; digit3<=MIN; end
      16'd725: begin digit0<=FIVE; digit1<=TWO; digit2<=SEVEN; digit3<=MIN; end
      16'd726: begin digit0<=SIX; digit1<=TWO; digit2<=SEVEN; digit3<=MIN; end
      16'd727: begin digit0<=SEVEN; digit1<=TWO; digit2<=SEVEN; digit3<=MIN; end
      16'd728: begin digit0<=EIGHT; digit1<=TWO; digit2<=SEVEN; digit3<=MIN; end
      16'd729: begin digit0<=NINE; digit1<=TWO; digit2<=SEVEN; digit3<=MIN; end
      16'd730: begin digit0<=ZERO; digit1<=THREE; digit2<=SEVEN; digit3<=MIN; end
      16'd731: begin digit0<=ONE; digit1<=THREE; digit2<=SEVEN; digit3<=MIN; end
      16'd732: begin digit0<=TWO; digit1<=THREE; digit2<=SEVEN; digit3<=MIN; end
      16'd733: begin digit0<=THREE; digit1<=THREE; digit2<=SEVEN; digit3<=MIN; end
      16'd734: begin digit0<=FOUR; digit1<=THREE; digit2<=SEVEN; digit3<=MIN; end
      16'd735: begin digit0<=FIVE; digit1<=THREE; digit2<=SEVEN; digit3<=MIN; end
      16'd736: begin digit0<=SIX; digit1<=THREE; digit2<=SEVEN; digit3<=MIN; end
      16'd737: begin digit0<=SEVEN; digit1<=THREE; digit2<=SEVEN; digit3<=MIN; end
      16'd738: begin digit0<=EIGHT; digit1<=THREE; digit2<=SEVEN; digit3<=MIN; end
      16'd739: begin digit0<=NINE; digit1<=THREE; digit2<=SEVEN; digit3<=MIN; end
      16'd740: begin digit0<=ZERO; digit1<=FOUR; digit2<=SEVEN; digit3<=MIN; end
      16'd741: begin digit0<=ONE; digit1<=FOUR; digit2<=SEVEN; digit3<=MIN; end
      16'd742: begin digit0<=TWO; digit1<=FOUR; digit2<=SEVEN; digit3<=MIN; end
      16'd743: begin digit0<=THREE; digit1<=FOUR; digit2<=SEVEN; digit3<=MIN; end
      16'd744: begin digit0<=FOUR; digit1<=FOUR; digit2<=SEVEN; digit3<=MIN; end
      16'd745: begin digit0<=FIVE; digit1<=FOUR; digit2<=SEVEN; digit3<=MIN; end
      16'd746: begin digit0<=SIX; digit1<=FOUR; digit2<=SEVEN; digit3<=MIN; end
      16'd747: begin digit0<=SEVEN; digit1<=FOUR; digit2<=SEVEN; digit3<=MIN; end
      16'd748: begin digit0<=EIGHT; digit1<=FOUR; digit2<=SEVEN; digit3<=MIN; end
      16'd749: begin digit0<=NINE; digit1<=FOUR; digit2<=SEVEN; digit3<=MIN; end
      16'd750: begin digit0<=ZERO; digit1<=FIVE; digit2<=SEVEN; digit3<=MIN; end
      16'd751: begin digit0<=ONE; digit1<=FIVE; digit2<=SEVEN; digit3<=MIN; end
      16'd752: begin digit0<=TWO; digit1<=FIVE; digit2<=SEVEN; digit3<=MIN; end
      16'd753: begin digit0<=THREE; digit1<=FIVE; digit2<=SEVEN; digit3<=MIN; end
      16'd754: begin digit0<=FOUR; digit1<=FIVE; digit2<=SEVEN; digit3<=MIN; end
      16'd755: begin digit0<=FIVE; digit1<=FIVE; digit2<=SEVEN; digit3<=MIN; end
      16'd756: begin digit0<=SIX; digit1<=FIVE; digit2<=SEVEN; digit3<=MIN; end
      16'd757: begin digit0<=SEVEN; digit1<=FIVE; digit2<=SEVEN; digit3<=MIN; end
      16'd758: begin digit0<=EIGHT; digit1<=FIVE; digit2<=SEVEN; digit3<=MIN; end
      16'd759: begin digit0<=NINE; digit1<=FIVE; digit2<=SEVEN; digit3<=MIN; end
      16'd760: begin digit0<=ZERO; digit1<=SIX; digit2<=SEVEN; digit3<=MIN; end
      16'd761: begin digit0<=ONE; digit1<=SIX; digit2<=SEVEN; digit3<=MIN; end
      16'd762: begin digit0<=TWO; digit1<=SIX; digit2<=SEVEN; digit3<=MIN; end
      16'd763: begin digit0<=THREE; digit1<=SIX; digit2<=SEVEN; digit3<=MIN; end
      16'd764: begin digit0<=FOUR; digit1<=SIX; digit2<=SEVEN; digit3<=MIN; end
      16'd765: begin digit0<=FIVE; digit1<=SIX; digit2<=SEVEN; digit3<=MIN; end
      16'd766: begin digit0<=SIX; digit1<=SIX; digit2<=SEVEN; digit3<=MIN; end
      16'd767: begin digit0<=SEVEN; digit1<=SIX; digit2<=SEVEN; digit3<=MIN; end
      16'd768: begin digit0<=EIGHT; digit1<=SIX; digit2<=SEVEN; digit3<=MIN; end
      16'd769: begin digit0<=NINE; digit1<=SIX; digit2<=SEVEN; digit3<=MIN; end
      16'd770: begin digit0<=ZERO; digit1<=SEVEN; digit2<=SEVEN; digit3<=MIN; end
      16'd771: begin digit0<=ONE; digit1<=SEVEN; digit2<=SEVEN; digit3<=MIN; end
      16'd772: begin digit0<=TWO; digit1<=SEVEN; digit2<=SEVEN; digit3<=MIN; end
      16'd773: begin digit0<=THREE; digit1<=SEVEN; digit2<=SEVEN; digit3<=MIN; end
      16'd774: begin digit0<=FOUR; digit1<=SEVEN; digit2<=SEVEN; digit3<=MIN; end
      16'd775: begin digit0<=FIVE; digit1<=SEVEN; digit2<=SEVEN; digit3<=MIN; end
      16'd776: begin digit0<=SIX; digit1<=SEVEN; digit2<=SEVEN; digit3<=MIN; end
      16'd777: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=SEVEN; digit3<=MIN; end
      16'd778: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=SEVEN; digit3<=MIN; end
      16'd779: begin digit0<=NINE; digit1<=SEVEN; digit2<=SEVEN; digit3<=MIN; end
      16'd780: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=MIN; end
      16'd781: begin digit0<=ONE; digit1<=EIGHT; digit2<=SEVEN; digit3<=MIN; end
      16'd782: begin digit0<=ZERO; digit1<=EIGHT; digit2<=SEVEN; digit3<=MIN; end
      16'd783: begin digit0<=THREE; digit1<=EIGHT; digit2<=SEVEN; digit3<=MIN; end
      16'd784: begin digit0<=FOUR; digit1<=EIGHT; digit2<=SEVEN; digit3<=MIN; end
      16'd785: begin digit0<=FIVE; digit1<=EIGHT; digit2<=SEVEN; digit3<=MIN; end
      16'd786: begin digit0<=SIX; digit1<=EIGHT; digit2<=SEVEN; digit3<=MIN; end
      16'd787: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=SEVEN; digit3<=MIN; end
      16'd788: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=SEVEN; digit3<=MIN; end
      16'd789: begin digit0<=NINE; digit1<=EIGHT; digit2<=SEVEN; digit3<=MIN; end
      16'd790: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=MIN; end
      16'd791: begin digit0<=ONE; digit1<=NINE; digit2<=SEVEN; digit3<=MIN; end
      16'd792: begin digit0<=ZERO; digit1<=NINE; digit2<=SEVEN; digit3<=MIN; end
      16'd793: begin digit0<=THREE; digit1<=NINE; digit2<=SEVEN; digit3<=MIN; end
      16'd794: begin digit0<=FOUR; digit1<=NINE; digit2<=SEVEN; digit3<=MIN; end
      16'd795: begin digit0<=FIVE; digit1<=NINE; digit2<=SEVEN; digit3<=MIN; end
      16'd796: begin digit0<=SIX; digit1<=NINE; digit2<=SEVEN; digit3<=MIN; end
      16'd797: begin digit0<=SEVEN; digit1<=NINE; digit2<=SEVEN; digit3<=MIN; end
      16'd798: begin digit0<=EIGHT; digit1<=NINE; digit2<=SEVEN; digit3<=MIN; end
      16'd799: begin digit0<=NINE; digit1<=NINE; digit2<=SEVEN; digit3<=MIN; end
	  16'd800: begin digit0<=ZERO; digit1<=ZERO; digit2<=EIGHT; digit3<=MIN; end
      16'd801: begin digit0<=ONE; digit1<=ZERO; digit2<=EIGHT; digit3<=MIN; end
      16'd802: begin digit0<=TWO; digit1<=ZERO; digit2<=EIGHT; digit3<=MIN; end
      16'd803: begin digit0<=THREE; digit1<=ZERO; digit2<=EIGHT; digit3<=MIN; end
      16'd804: begin digit0<=FOUR; digit1<=ZERO; digit2<=EIGHT; digit3<=MIN; end
      16'd805: begin digit0<=FIVE; digit1<=ZERO; digit2<=EIGHT; digit3<=MIN; end
      16'd806: begin digit0<=SIX; digit1<=ZERO; digit2<=EIGHT; digit3<=MIN; end
      16'd807: begin digit0<=SEVEN; digit1<=ZERO; digit2<=EIGHT; digit3<=MIN; end
      16'd808: begin digit0<=EIGHT; digit1<=ZERO; digit2<=EIGHT; digit3<=MIN; end
      16'd809: begin digit0<=NINE; digit1<=ZERO; digit2<=EIGHT; digit3<=MIN; end
      16'd810: begin digit0<=ZERO; digit1<=ONE; digit2<=EIGHT; digit3<=MIN; end
      16'd811: begin digit0<=ONE; digit1<=ONE; digit2<=EIGHT; digit3<=MIN; end
      16'd812: begin digit0<=TWO; digit1<=ONE; digit2<=EIGHT; digit3<=MIN; end
      16'd813: begin digit0<=THREE; digit1<=ONE; digit2<=EIGHT; digit3<=MIN; end
      16'd814: begin digit0<=FOUR; digit1<=ONE; digit2<=EIGHT; digit3<=MIN; end
      16'd815: begin digit0<=FIVE; digit1<=ONE; digit2<=EIGHT; digit3<=MIN; end
      16'd816: begin digit0<=SIX; digit1<=ONE; digit2<=EIGHT; digit3<=MIN; end
      16'd817: begin digit0<=SEVEN; digit1<=ONE; digit2<=EIGHT; digit3<=MIN; end
      16'd818: begin digit0<=EIGHT; digit1<=ONE; digit2<=EIGHT; digit3<=MIN; end
      16'd819: begin digit0<=NINE; digit1<=ONE; digit2<=EIGHT; digit3<=MIN; end
      16'd820: begin digit0<=ZERO; digit1<=TWO; digit2<=EIGHT; digit3<=MIN; end
      16'd821: begin digit0<=ONE; digit1<=TWO; digit2<=EIGHT; digit3<=MIN; end
      16'd822: begin digit0<=TWO; digit1<=TWO; digit2<=EIGHT; digit3<=MIN; end
      16'd823: begin digit0<=THREE; digit1<=TWO; digit2<=EIGHT; digit3<=MIN; end
      16'd824: begin digit0<=FOUR; digit1<=TWO; digit2<=EIGHT; digit3<=MIN; end
      16'd825: begin digit0<=FIVE; digit1<=TWO; digit2<=EIGHT; digit3<=MIN; end
      16'd826: begin digit0<=SIX; digit1<=TWO; digit2<=EIGHT; digit3<=MIN; end
      16'd827: begin digit0<=SEVEN; digit1<=TWO; digit2<=EIGHT; digit3<=MIN; end
      16'd828: begin digit0<=EIGHT; digit1<=TWO; digit2<=EIGHT; digit3<=MIN; end
      16'd829: begin digit0<=NINE; digit1<=TWO; digit2<=EIGHT; digit3<=MIN; end
      16'd830: begin digit0<=ZERO; digit1<=THREE; digit2<=EIGHT; digit3<=MIN; end
      16'd831: begin digit0<=ONE; digit1<=THREE; digit2<=EIGHT; digit3<=MIN; end
      16'd832: begin digit0<=TWO; digit1<=THREE; digit2<=EIGHT; digit3<=MIN; end
      16'd833: begin digit0<=THREE; digit1<=THREE; digit2<=EIGHT; digit3<=MIN; end
      16'd834: begin digit0<=FOUR; digit1<=THREE; digit2<=EIGHT; digit3<=MIN; end
      16'd835: begin digit0<=FIVE; digit1<=THREE; digit2<=EIGHT; digit3<=MIN; end
      16'd836: begin digit0<=SIX; digit1<=THREE; digit2<=EIGHT; digit3<=MIN; end
      16'd837: begin digit0<=SEVEN; digit1<=THREE; digit2<=EIGHT; digit3<=MIN; end
      16'd838: begin digit0<=EIGHT; digit1<=THREE; digit2<=EIGHT; digit3<=MIN; end
      16'd839: begin digit0<=NINE; digit1<=THREE; digit2<=EIGHT; digit3<=MIN; end
      16'd840: begin digit0<=ZERO; digit1<=FOUR; digit2<=EIGHT; digit3<=MIN; end
      16'd841: begin digit0<=ONE; digit1<=FOUR; digit2<=EIGHT; digit3<=MIN; end
      16'd842: begin digit0<=TWO; digit1<=FOUR; digit2<=EIGHT; digit3<=MIN; end
      16'd843: begin digit0<=THREE; digit1<=FOUR; digit2<=EIGHT; digit3<=MIN; end
      16'd844: begin digit0<=FOUR; digit1<=FOUR; digit2<=EIGHT; digit3<=MIN; end
      16'd845: begin digit0<=FIVE; digit1<=FOUR; digit2<=EIGHT; digit3<=MIN; end
      16'd846: begin digit0<=SIX; digit1<=FOUR; digit2<=EIGHT; digit3<=MIN; end
      16'd847: begin digit0<=SEVEN; digit1<=FOUR; digit2<=EIGHT; digit3<=MIN; end
      16'd848: begin digit0<=EIGHT; digit1<=FOUR; digit2<=EIGHT; digit3<=MIN; end
      16'd849: begin digit0<=NINE; digit1<=FOUR; digit2<=EIGHT; digit3<=MIN; end
      16'd850: begin digit0<=ZERO; digit1<=FIVE; digit2<=EIGHT; digit3<=MIN; end
      16'd851: begin digit0<=ONE; digit1<=FIVE; digit2<=EIGHT; digit3<=MIN; end
      16'd852: begin digit0<=TWO; digit1<=FIVE; digit2<=EIGHT; digit3<=MIN; end
      16'd853: begin digit0<=THREE; digit1<=FIVE; digit2<=EIGHT; digit3<=MIN; end
      16'd854: begin digit0<=FOUR; digit1<=FIVE; digit2<=EIGHT; digit3<=MIN; end
      16'd855: begin digit0<=FIVE; digit1<=FIVE; digit2<=EIGHT; digit3<=MIN; end
      16'd856: begin digit0<=SIX; digit1<=FIVE; digit2<=EIGHT; digit3<=MIN; end
      16'd857: begin digit0<=SEVEN; digit1<=FIVE; digit2<=EIGHT; digit3<=MIN; end
      16'd858: begin digit0<=EIGHT; digit1<=FIVE; digit2<=EIGHT; digit3<=MIN; end
      16'd859: begin digit0<=NINE; digit1<=FIVE; digit2<=EIGHT; digit3<=MIN; end
      16'd860: begin digit0<=ZERO; digit1<=SIX; digit2<=EIGHT; digit3<=MIN; end
      16'd861: begin digit0<=ONE; digit1<=SIX; digit2<=EIGHT; digit3<=MIN; end
      16'd862: begin digit0<=TWO; digit1<=SIX; digit2<=EIGHT; digit3<=MIN; end
      16'd863: begin digit0<=THREE; digit1<=SIX; digit2<=EIGHT; digit3<=MIN; end
      16'd864: begin digit0<=FOUR; digit1<=SIX; digit2<=EIGHT; digit3<=MIN; end
      16'd865: begin digit0<=FIVE; digit1<=SIX; digit2<=EIGHT; digit3<=MIN; end
      16'd866: begin digit0<=SIX; digit1<=SIX; digit2<=EIGHT; digit3<=MIN; end
      16'd867: begin digit0<=SEVEN; digit1<=SIX; digit2<=EIGHT; digit3<=MIN; end
      16'd868: begin digit0<=EIGHT; digit1<=SIX; digit2<=EIGHT; digit3<=MIN; end
      16'd869: begin digit0<=NINE; digit1<=SIX; digit2<=EIGHT; digit3<=MIN; end
      16'd870: begin digit0<=ZERO; digit1<=SEVEN; digit2<=EIGHT; digit3<=MIN; end
      16'd871: begin digit0<=ONE; digit1<=SEVEN; digit2<=EIGHT; digit3<=MIN; end
      16'd872: begin digit0<=TWO; digit1<=SEVEN; digit2<=EIGHT; digit3<=MIN; end
      16'd873: begin digit0<=THREE; digit1<=SEVEN; digit2<=EIGHT; digit3<=MIN; end
      16'd874: begin digit0<=FOUR; digit1<=SEVEN; digit2<=EIGHT; digit3<=MIN; end
      16'd875: begin digit0<=FIVE; digit1<=SEVEN; digit2<=EIGHT; digit3<=MIN; end
      16'd876: begin digit0<=SIX; digit1<=SEVEN; digit2<=EIGHT; digit3<=MIN; end
      16'd877: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=EIGHT; digit3<=MIN; end
      16'd878: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=EIGHT; digit3<=MIN; end
      16'd879: begin digit0<=NINE; digit1<=SEVEN; digit2<=EIGHT; digit3<=MIN; end
      16'd880: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=MIN; end
      16'd881: begin digit0<=ONE; digit1<=EIGHT; digit2<=EIGHT; digit3<=MIN; end
      16'd882: begin digit0<=ZERO; digit1<=EIGHT; digit2<=EIGHT; digit3<=MIN; end
      16'd883: begin digit0<=THREE; digit1<=EIGHT; digit2<=EIGHT; digit3<=MIN; end
      16'd884: begin digit0<=FOUR; digit1<=EIGHT; digit2<=EIGHT; digit3<=MIN; end
      16'd885: begin digit0<=FIVE; digit1<=EIGHT; digit2<=EIGHT; digit3<=MIN; end
      16'd886: begin digit0<=SIX; digit1<=EIGHT; digit2<=EIGHT; digit3<=MIN; end
      16'd887: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=EIGHT; digit3<=MIN; end
      16'd888: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=EIGHT; digit3<=MIN; end
      16'd889: begin digit0<=NINE; digit1<=EIGHT; digit2<=EIGHT; digit3<=MIN; end
      16'd890: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=MIN; end
      16'd891: begin digit0<=ONE; digit1<=NINE; digit2<=EIGHT; digit3<=MIN; end
      16'd892: begin digit0<=ZERO; digit1<=NINE; digit2<=EIGHT; digit3<=MIN; end
      16'd893: begin digit0<=THREE; digit1<=NINE; digit2<=EIGHT; digit3<=MIN; end
      16'd894: begin digit0<=FOUR; digit1<=NINE; digit2<=EIGHT; digit3<=MIN; end
      16'd895: begin digit0<=FIVE; digit1<=NINE; digit2<=EIGHT; digit3<=MIN; end
      16'd896: begin digit0<=SIX; digit1<=NINE; digit2<=EIGHT; digit3<=MIN; end
      16'd897: begin digit0<=SEVEN; digit1<=NINE; digit2<=EIGHT; digit3<=MIN; end
      16'd898: begin digit0<=EIGHT; digit1<=NINE; digit2<=EIGHT; digit3<=MIN; end
      16'd899: begin digit0<=NINE; digit1<=NINE; digit2<=EIGHT; digit3<=MIN; end
	  16'd900: begin digit0<=ZERO; digit1<=ZERO; digit2<=NINE; digit3<=MIN; end
      16'd901: begin digit0<=ONE; digit1<=ZERO; digit2<=NINE; digit3<=MIN; end
      16'd902: begin digit0<=TWO; digit1<=ZERO; digit2<=NINE; digit3<=MIN; end
      16'd903: begin digit0<=THREE; digit1<=ZERO; digit2<=NINE; digit3<=MIN; end
      16'd904: begin digit0<=FOUR; digit1<=ZERO; digit2<=NINE; digit3<=MIN; end
      16'd905: begin digit0<=FIVE; digit1<=ZERO; digit2<=NINE; digit3<=MIN; end
      16'd906: begin digit0<=SIX; digit1<=ZERO; digit2<=NINE; digit3<=MIN; end
      16'd907: begin digit0<=SEVEN; digit1<=ZERO; digit2<=NINE; digit3<=MIN; end
      16'd908: begin digit0<=EIGHT; digit1<=ZERO; digit2<=NINE; digit3<=MIN; end
      16'd909: begin digit0<=NINE; digit1<=ZERO; digit2<=NINE; digit3<=MIN; end
      16'd910: begin digit0<=ZERO; digit1<=ONE; digit2<=NINE; digit3<=MIN; end
      16'd911: begin digit0<=ONE; digit1<=ONE; digit2<=NINE; digit3<=MIN; end
      16'd912: begin digit0<=TWO; digit1<=ONE; digit2<=NINE; digit3<=MIN; end
      16'd913: begin digit0<=THREE; digit1<=ONE; digit2<=NINE; digit3<=MIN; end
      16'd914: begin digit0<=FOUR; digit1<=ONE; digit2<=NINE; digit3<=MIN; end
      16'd915: begin digit0<=FIVE; digit1<=ONE; digit2<=NINE; digit3<=MIN; end
      16'd916: begin digit0<=SIX; digit1<=ONE; digit2<=NINE; digit3<=MIN; end
      16'd917: begin digit0<=SEVEN; digit1<=ONE; digit2<=NINE; digit3<=MIN; end
      16'd918: begin digit0<=EIGHT; digit1<=ONE; digit2<=NINE; digit3<=MIN; end
      16'd919: begin digit0<=NINE; digit1<=ONE; digit2<=NINE; digit3<=MIN; end
      16'd920: begin digit0<=ZERO; digit1<=TWO; digit2<=NINE; digit3<=MIN; end
      16'd921: begin digit0<=ONE; digit1<=TWO; digit2<=NINE; digit3<=MIN; end
      16'd922: begin digit0<=TWO; digit1<=TWO; digit2<=NINE; digit3<=MIN; end
      16'd923: begin digit0<=THREE; digit1<=TWO; digit2<=NINE; digit3<=MIN; end
      16'd924: begin digit0<=FOUR; digit1<=TWO; digit2<=NINE; digit3<=MIN; end
      16'd925: begin digit0<=FIVE; digit1<=TWO; digit2<=NINE; digit3<=MIN; end
      16'd926: begin digit0<=SIX; digit1<=TWO; digit2<=NINE; digit3<=MIN; end
      16'd927: begin digit0<=SEVEN; digit1<=TWO; digit2<=NINE; digit3<=MIN; end
      16'd928: begin digit0<=EIGHT; digit1<=TWO; digit2<=NINE; digit3<=MIN; end
      16'd929: begin digit0<=NINE; digit1<=TWO; digit2<=NINE; digit3<=MIN; end
      16'd930: begin digit0<=ZERO; digit1<=THREE; digit2<=NINE; digit3<=MIN; end
      16'd931: begin digit0<=ONE; digit1<=THREE; digit2<=NINE; digit3<=MIN; end
      16'd932: begin digit0<=TWO; digit1<=THREE; digit2<=NINE; digit3<=MIN; end
      16'd933: begin digit0<=THREE; digit1<=THREE; digit2<=NINE; digit3<=MIN; end
      16'd934: begin digit0<=FOUR; digit1<=THREE; digit2<=NINE; digit3<=MIN; end
      16'd935: begin digit0<=FIVE; digit1<=THREE; digit2<=NINE; digit3<=MIN; end
      16'd936: begin digit0<=SIX; digit1<=THREE; digit2<=NINE; digit3<=MIN; end
      16'd937: begin digit0<=SEVEN; digit1<=THREE; digit2<=NINE; digit3<=MIN; end
      16'd938: begin digit0<=EIGHT; digit1<=THREE; digit2<=NINE; digit3<=MIN; end
      16'd939: begin digit0<=NINE; digit1<=THREE; digit2<=NINE; digit3<=MIN; end
      16'd940: begin digit0<=ZERO; digit1<=FOUR; digit2<=NINE; digit3<=MIN; end
      16'd941: begin digit0<=ONE; digit1<=FOUR; digit2<=NINE; digit3<=MIN; end
      16'd942: begin digit0<=TWO; digit1<=FOUR; digit2<=NINE; digit3<=MIN; end
      16'd943: begin digit0<=THREE; digit1<=FOUR; digit2<=NINE; digit3<=MIN; end
      16'd944: begin digit0<=FOUR; digit1<=FOUR; digit2<=NINE; digit3<=MIN; end
      16'd945: begin digit0<=FIVE; digit1<=FOUR; digit2<=NINE; digit3<=MIN; end
      16'd946: begin digit0<=SIX; digit1<=FOUR; digit2<=NINE; digit3<=MIN; end
      16'd947: begin digit0<=SEVEN; digit1<=FOUR; digit2<=NINE; digit3<=MIN; end
      16'd948: begin digit0<=EIGHT; digit1<=FOUR; digit2<=NINE; digit3<=MIN; end
      16'd949: begin digit0<=NINE; digit1<=FOUR; digit2<=NINE; digit3<=MIN; end
      16'd950: begin digit0<=ZERO; digit1<=FIVE; digit2<=NINE; digit3<=MIN; end
      16'd951: begin digit0<=ONE; digit1<=FIVE; digit2<=NINE; digit3<=MIN; end
      16'd952: begin digit0<=TWO; digit1<=FIVE; digit2<=NINE; digit3<=MIN; end
      16'd953: begin digit0<=THREE; digit1<=FIVE; digit2<=NINE; digit3<=MIN; end
      16'd954: begin digit0<=FOUR; digit1<=FIVE; digit2<=NINE; digit3<=MIN; end
      16'd955: begin digit0<=FIVE; digit1<=FIVE; digit2<=NINE; digit3<=MIN; end
      16'd956: begin digit0<=SIX; digit1<=FIVE; digit2<=NINE; digit3<=MIN; end
      16'd957: begin digit0<=SEVEN; digit1<=FIVE; digit2<=NINE; digit3<=MIN; end
      16'd958: begin digit0<=EIGHT; digit1<=FIVE; digit2<=NINE; digit3<=MIN; end
      16'd959: begin digit0<=NINE; digit1<=FIVE; digit2<=NINE; digit3<=MIN; end
      16'd960: begin digit0<=ZERO; digit1<=SIX; digit2<=NINE; digit3<=MIN; end
      16'd961: begin digit0<=ONE; digit1<=SIX; digit2<=NINE; digit3<=MIN; end
      16'd962: begin digit0<=TWO; digit1<=SIX; digit2<=NINE; digit3<=MIN; end
      16'd963: begin digit0<=THREE; digit1<=SIX; digit2<=NINE; digit3<=MIN; end
      16'd964: begin digit0<=FOUR; digit1<=SIX; digit2<=NINE; digit3<=MIN; end
      16'd965: begin digit0<=FIVE; digit1<=SIX; digit2<=NINE; digit3<=MIN; end
      16'd966: begin digit0<=SIX; digit1<=SIX; digit2<=NINE; digit3<=MIN; end
      16'd967: begin digit0<=SEVEN; digit1<=SIX; digit2<=NINE; digit3<=MIN; end
      16'd968: begin digit0<=EIGHT; digit1<=SIX; digit2<=NINE; digit3<=MIN; end
      16'd969: begin digit0<=NINE; digit1<=SIX; digit2<=NINE; digit3<=MIN; end
      16'd970: begin digit0<=ZERO; digit1<=SEVEN; digit2<=NINE; digit3<=MIN; end
      16'd971: begin digit0<=ONE; digit1<=SEVEN; digit2<=NINE; digit3<=MIN; end
      16'd972: begin digit0<=TWO; digit1<=SEVEN; digit2<=NINE; digit3<=MIN; end
      16'd973: begin digit0<=THREE; digit1<=SEVEN; digit2<=NINE; digit3<=MIN; end
      16'd974: begin digit0<=FOUR; digit1<=SEVEN; digit2<=NINE; digit3<=MIN; end
      16'd975: begin digit0<=FIVE; digit1<=SEVEN; digit2<=NINE; digit3<=MIN; end
      16'd976: begin digit0<=SIX; digit1<=SEVEN; digit2<=NINE; digit3<=MIN; end
      16'd977: begin digit0<=SEVEN; digit1<=SEVEN; digit2<=NINE; digit3<=MIN; end
      16'd978: begin digit0<=EIGHT; digit1<=SEVEN; digit2<=NINE; digit3<=MIN; end
      16'd979: begin digit0<=NINE; digit1<=SEVEN; digit2<=NINE; digit3<=MIN; end
      16'd980: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=MIN; end
      16'd981: begin digit0<=ONE; digit1<=EIGHT; digit2<=NINE; digit3<=MIN; end
      16'd982: begin digit0<=ZERO; digit1<=EIGHT; digit2<=NINE; digit3<=MIN; end
      16'd983: begin digit0<=THREE; digit1<=EIGHT; digit2<=NINE; digit3<=MIN; end
      16'd984: begin digit0<=FOUR; digit1<=EIGHT; digit2<=NINE; digit3<=MIN; end
      16'd985: begin digit0<=FIVE; digit1<=EIGHT; digit2<=NINE; digit3<=MIN; end
      16'd986: begin digit0<=SIX; digit1<=EIGHT; digit2<=NINE; digit3<=MIN; end
      16'd987: begin digit0<=SEVEN; digit1<=EIGHT; digit2<=NINE; digit3<=MIN; end
      16'd988: begin digit0<=EIGHT; digit1<=EIGHT; digit2<=NINE; digit3<=MIN; end
      16'd989: begin digit0<=NINE; digit1<=EIGHT; digit2<=NINE; digit3<=MIN; end
      16'd990: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=MIN; end
      16'd991: begin digit0<=ONE; digit1<=NINE; digit2<=NINE; digit3<=MIN; end
      16'd992: begin digit0<=ZERO; digit1<=NINE; digit2<=NINE; digit3<=MIN; end
      16'd993: begin digit0<=THREE; digit1<=NINE; digit2<=NINE; digit3<=MIN; end
      16'd994: begin digit0<=FOUR; digit1<=NINE; digit2<=NINE; digit3<=MIN; end
      16'd995: begin digit0<=FIVE; digit1<=NINE; digit2<=NINE; digit3<=MIN; end
      16'd996: begin digit0<=SIX; digit1<=NINE; digit2<=NINE; digit3<=MIN; end
      16'd997: begin digit0<=SEVEN; digit1<=NINE; digit2<=NINE; digit3<=MIN; end
      16'd998: begin digit0<=EIGHT; digit1<=NINE; digit2<=NINE; digit3<=MIN; end
      16'd999: begin digit0<=NINE; digit1<=NINE; digit2<=NINE; digit3<=MIN; end
      default: begin digit0<=EMPTY; digit1<=EMPTY; digit2<=EMPTY; digit3<=EMPTY; end
    endcase
  else 
      begin
      digit0<=EMPTY;
      digit1<=EMPTY;
	  digit2<=EMPTY;
	  digit3<=EMPTY;
      end
end
endmodule
